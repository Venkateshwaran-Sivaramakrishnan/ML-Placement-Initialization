module aes_cipher_top (clk,
    done,
    ld,
    rst,
    key,
    text_in,
    text_out);
 input clk;
 output done;
 input ld;
 input rst;
 input [127:0] key;
 input [127:0] text_in;
 output [127:0] text_out;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire net836;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire net188;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire net870;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire net806;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire net126;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire net162;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire net724;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire net203;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire net3;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire net733;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire net200;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire net202;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire net156;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire net2;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire net154;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire net157;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire net155;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire net195;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire net196;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire net197;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire net13;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire net161;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire net97;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire net1113;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire net32;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire net6;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire net159;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire net958;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire net106;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire net14;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire net108;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire net568;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire net628;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire net1199;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire net1225;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire net1166;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire net828;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire _06406_;
 wire _06407_;
 wire _06408_;
 wire _06409_;
 wire _06410_;
 wire _06411_;
 wire _06412_;
 wire _06413_;
 wire _06414_;
 wire _06415_;
 wire _06416_;
 wire _06417_;
 wire _06418_;
 wire _06419_;
 wire _06420_;
 wire _06421_;
 wire _06422_;
 wire _06423_;
 wire _06424_;
 wire _06425_;
 wire _06426_;
 wire _06427_;
 wire _06428_;
 wire _06429_;
 wire _06430_;
 wire _06431_;
 wire _06432_;
 wire _06433_;
 wire _06434_;
 wire _06435_;
 wire _06436_;
 wire _06437_;
 wire _06438_;
 wire _06439_;
 wire _06440_;
 wire _06441_;
 wire _06442_;
 wire _06443_;
 wire _06444_;
 wire _06445_;
 wire _06446_;
 wire _06447_;
 wire _06448_;
 wire _06449_;
 wire _06450_;
 wire _06451_;
 wire _06452_;
 wire _06453_;
 wire _06454_;
 wire _06455_;
 wire _06456_;
 wire _06457_;
 wire _06458_;
 wire _06459_;
 wire _06460_;
 wire _06461_;
 wire _06462_;
 wire _06463_;
 wire _06464_;
 wire _06465_;
 wire _06466_;
 wire _06467_;
 wire _06468_;
 wire _06469_;
 wire _06470_;
 wire net1048;
 wire _06472_;
 wire _06473_;
 wire _06474_;
 wire _06475_;
 wire _06476_;
 wire _06477_;
 wire _06478_;
 wire _06479_;
 wire _06480_;
 wire _06481_;
 wire _06482_;
 wire _06483_;
 wire _06484_;
 wire _06485_;
 wire _06486_;
 wire _06487_;
 wire _06488_;
 wire _06489_;
 wire _06490_;
 wire _06491_;
 wire _06492_;
 wire _06493_;
 wire _06494_;
 wire _06495_;
 wire _06496_;
 wire _06497_;
 wire _06498_;
 wire _06499_;
 wire _06500_;
 wire _06501_;
 wire _06502_;
 wire _06503_;
 wire _06504_;
 wire _06505_;
 wire _06506_;
 wire _06507_;
 wire _06508_;
 wire _06509_;
 wire _06510_;
 wire _06511_;
 wire _06512_;
 wire _06513_;
 wire _06514_;
 wire _06515_;
 wire _06516_;
 wire _06517_;
 wire _06518_;
 wire _06519_;
 wire _06520_;
 wire _06521_;
 wire _06522_;
 wire _06523_;
 wire _06524_;
 wire _06525_;
 wire _06526_;
 wire _06527_;
 wire _06528_;
 wire _06529_;
 wire _06530_;
 wire _06531_;
 wire _06532_;
 wire _06533_;
 wire _06534_;
 wire _06535_;
 wire _06536_;
 wire _06537_;
 wire _06538_;
 wire _06539_;
 wire _06540_;
 wire _06541_;
 wire _06542_;
 wire _06543_;
 wire _06544_;
 wire _06545_;
 wire _06546_;
 wire _06547_;
 wire _06548_;
 wire _06549_;
 wire _06550_;
 wire _06551_;
 wire _06552_;
 wire _06553_;
 wire _06554_;
 wire _06555_;
 wire _06556_;
 wire _06557_;
 wire _06558_;
 wire _06559_;
 wire _06560_;
 wire _06561_;
 wire _06562_;
 wire _06563_;
 wire _06564_;
 wire _06565_;
 wire _06566_;
 wire _06567_;
 wire _06568_;
 wire _06569_;
 wire _06570_;
 wire _06571_;
 wire _06572_;
 wire _06573_;
 wire _06574_;
 wire _06575_;
 wire _06576_;
 wire _06577_;
 wire _06578_;
 wire _06579_;
 wire _06580_;
 wire _06581_;
 wire _06582_;
 wire _06583_;
 wire _06584_;
 wire _06585_;
 wire _06586_;
 wire _06587_;
 wire _06588_;
 wire _06589_;
 wire _06590_;
 wire _06591_;
 wire _06592_;
 wire _06593_;
 wire _06594_;
 wire _06595_;
 wire _06596_;
 wire _06597_;
 wire _06598_;
 wire _06599_;
 wire _06600_;
 wire _06601_;
 wire net786;
 wire _06603_;
 wire _06604_;
 wire net782;
 wire _06606_;
 wire _06607_;
 wire _06608_;
 wire _06609_;
 wire _06610_;
 wire _06611_;
 wire _06612_;
 wire _06613_;
 wire _06614_;
 wire _06615_;
 wire _06616_;
 wire _06617_;
 wire _06618_;
 wire _06619_;
 wire _06620_;
 wire net795;
 wire net1087;
 wire _06623_;
 wire _06624_;
 wire _06625_;
 wire _06626_;
 wire _06627_;
 wire _06628_;
 wire _06629_;
 wire _06630_;
 wire _06631_;
 wire _06632_;
 wire _06633_;
 wire _06634_;
 wire _06635_;
 wire _06636_;
 wire _06637_;
 wire _06638_;
 wire _06639_;
 wire _06640_;
 wire _06641_;
 wire _06642_;
 wire _06643_;
 wire _06644_;
 wire _06645_;
 wire _06646_;
 wire _06647_;
 wire _06648_;
 wire _06649_;
 wire _06650_;
 wire _06651_;
 wire _06652_;
 wire _06653_;
 wire _06654_;
 wire _06655_;
 wire _06656_;
 wire _06657_;
 wire _06658_;
 wire _06659_;
 wire _06660_;
 wire _06661_;
 wire _06662_;
 wire _06663_;
 wire _06664_;
 wire _06665_;
 wire _06666_;
 wire _06667_;
 wire _06668_;
 wire _06669_;
 wire _06670_;
 wire _06671_;
 wire _06672_;
 wire _06673_;
 wire _06674_;
 wire _06675_;
 wire _06676_;
 wire _06677_;
 wire _06678_;
 wire _06679_;
 wire _06680_;
 wire _06681_;
 wire _06682_;
 wire _06683_;
 wire _06684_;
 wire _06685_;
 wire _06686_;
 wire _06687_;
 wire _06688_;
 wire _06689_;
 wire _06690_;
 wire _06691_;
 wire _06692_;
 wire _06693_;
 wire _06694_;
 wire _06695_;
 wire _06696_;
 wire _06697_;
 wire _06698_;
 wire _06699_;
 wire _06700_;
 wire _06701_;
 wire _06702_;
 wire _06703_;
 wire _06704_;
 wire _06705_;
 wire _06706_;
 wire _06707_;
 wire _06708_;
 wire _06709_;
 wire _06710_;
 wire _06711_;
 wire _06712_;
 wire _06713_;
 wire _06714_;
 wire _06715_;
 wire _06716_;
 wire _06717_;
 wire _06718_;
 wire _06719_;
 wire _06720_;
 wire _06721_;
 wire _06722_;
 wire _06723_;
 wire _06724_;
 wire _06725_;
 wire _06726_;
 wire _06727_;
 wire _06728_;
 wire _06729_;
 wire _06730_;
 wire _06731_;
 wire _06732_;
 wire _06733_;
 wire _06734_;
 wire _06735_;
 wire _06736_;
 wire _06737_;
 wire _06738_;
 wire _06739_;
 wire _06740_;
 wire _06741_;
 wire _06742_;
 wire _06743_;
 wire _06744_;
 wire _06745_;
 wire _06746_;
 wire _06747_;
 wire _06748_;
 wire _06749_;
 wire _06750_;
 wire _06751_;
 wire _06752_;
 wire _06753_;
 wire _06754_;
 wire _06755_;
 wire _06756_;
 wire _06757_;
 wire _06758_;
 wire _06759_;
 wire _06760_;
 wire _06761_;
 wire _06762_;
 wire _06763_;
 wire _06764_;
 wire _06765_;
 wire _06766_;
 wire _06767_;
 wire _06768_;
 wire _06769_;
 wire _06770_;
 wire _06771_;
 wire _06772_;
 wire _06773_;
 wire _06774_;
 wire _06775_;
 wire _06776_;
 wire _06777_;
 wire _06778_;
 wire _06779_;
 wire _06780_;
 wire _06781_;
 wire _06782_;
 wire _06783_;
 wire _06784_;
 wire _06785_;
 wire _06786_;
 wire _06787_;
 wire _06788_;
 wire _06789_;
 wire _06790_;
 wire _06791_;
 wire _06792_;
 wire _06793_;
 wire _06794_;
 wire _06795_;
 wire _06796_;
 wire _06797_;
 wire _06798_;
 wire _06799_;
 wire _06800_;
 wire _06801_;
 wire _06802_;
 wire _06803_;
 wire _06804_;
 wire _06805_;
 wire _06806_;
 wire _06807_;
 wire _06808_;
 wire _06809_;
 wire _06810_;
 wire _06811_;
 wire _06812_;
 wire _06813_;
 wire _06814_;
 wire _06815_;
 wire _06816_;
 wire _06817_;
 wire _06818_;
 wire _06819_;
 wire _06820_;
 wire _06821_;
 wire _06822_;
 wire _06823_;
 wire _06824_;
 wire _06825_;
 wire _06826_;
 wire _06827_;
 wire _06828_;
 wire _06829_;
 wire _06830_;
 wire _06831_;
 wire _06832_;
 wire _06833_;
 wire _06834_;
 wire _06835_;
 wire _06836_;
 wire _06837_;
 wire _06838_;
 wire _06839_;
 wire _06840_;
 wire _06841_;
 wire _06842_;
 wire _06843_;
 wire _06844_;
 wire _06845_;
 wire _06846_;
 wire _06847_;
 wire _06848_;
 wire _06849_;
 wire _06850_;
 wire _06851_;
 wire _06852_;
 wire _06853_;
 wire _06854_;
 wire _06855_;
 wire _06856_;
 wire _06857_;
 wire _06858_;
 wire _06859_;
 wire _06860_;
 wire _06861_;
 wire _06862_;
 wire _06863_;
 wire _06864_;
 wire _06865_;
 wire _06866_;
 wire _06867_;
 wire _06868_;
 wire _06869_;
 wire _06870_;
 wire net1028;
 wire _06872_;
 wire _06873_;
 wire _06874_;
 wire net42;
 wire _06876_;
 wire _06877_;
 wire _06878_;
 wire _06879_;
 wire _06880_;
 wire _06881_;
 wire _06882_;
 wire _06883_;
 wire _06884_;
 wire _06885_;
 wire _06886_;
 wire _06887_;
 wire net1204;
 wire _06889_;
 wire _06890_;
 wire _06891_;
 wire _06892_;
 wire _06893_;
 wire _06894_;
 wire _06895_;
 wire _06896_;
 wire _06897_;
 wire _06898_;
 wire _06899_;
 wire _06900_;
 wire _06901_;
 wire _06902_;
 wire _06903_;
 wire _06904_;
 wire _06905_;
 wire net64;
 wire _06907_;
 wire _06908_;
 wire net94;
 wire _06910_;
 wire _06911_;
 wire _06912_;
 wire _06913_;
 wire _06914_;
 wire _06915_;
 wire _06916_;
 wire _06917_;
 wire _06918_;
 wire _06919_;
 wire _06920_;
 wire _06921_;
 wire _06922_;
 wire net930;
 wire _06924_;
 wire _06925_;
 wire _06926_;
 wire _06927_;
 wire _06928_;
 wire _06929_;
 wire _06930_;
 wire _06931_;
 wire _06932_;
 wire _06933_;
 wire _06934_;
 wire _06935_;
 wire _06936_;
 wire _06937_;
 wire _06938_;
 wire net1193;
 wire _06940_;
 wire _06941_;
 wire _06942_;
 wire _06943_;
 wire _06944_;
 wire _06945_;
 wire _06946_;
 wire _06947_;
 wire _06948_;
 wire _06949_;
 wire _06950_;
 wire _06951_;
 wire _06952_;
 wire _06953_;
 wire _06954_;
 wire _06955_;
 wire _06956_;
 wire _06957_;
 wire _06958_;
 wire _06959_;
 wire _06960_;
 wire _06961_;
 wire _06962_;
 wire _06963_;
 wire _06964_;
 wire _06965_;
 wire _06966_;
 wire _06967_;
 wire _06968_;
 wire _06969_;
 wire _06970_;
 wire _06971_;
 wire _06972_;
 wire _06973_;
 wire _06974_;
 wire _06975_;
 wire _06976_;
 wire _06977_;
 wire _06978_;
 wire _06979_;
 wire _06980_;
 wire _06981_;
 wire _06982_;
 wire _06983_;
 wire _06984_;
 wire _06985_;
 wire _06986_;
 wire _06987_;
 wire _06988_;
 wire _06989_;
 wire _06990_;
 wire _06991_;
 wire _06992_;
 wire _06993_;
 wire _06994_;
 wire _06995_;
 wire _06996_;
 wire _06997_;
 wire _06998_;
 wire _06999_;
 wire _07000_;
 wire _07001_;
 wire _07002_;
 wire _07003_;
 wire _07004_;
 wire _07005_;
 wire _07006_;
 wire _07007_;
 wire _07008_;
 wire _07009_;
 wire _07010_;
 wire _07011_;
 wire _07012_;
 wire _07013_;
 wire _07014_;
 wire _07015_;
 wire _07016_;
 wire _07017_;
 wire _07018_;
 wire _07019_;
 wire _07020_;
 wire _07021_;
 wire _07022_;
 wire _07023_;
 wire _07024_;
 wire _07025_;
 wire _07026_;
 wire _07027_;
 wire _07028_;
 wire _07029_;
 wire _07030_;
 wire _07031_;
 wire _07032_;
 wire _07033_;
 wire _07034_;
 wire _07035_;
 wire _07036_;
 wire _07037_;
 wire _07038_;
 wire _07039_;
 wire _07040_;
 wire _07041_;
 wire _07042_;
 wire _07043_;
 wire _07044_;
 wire _07045_;
 wire _07046_;
 wire _07047_;
 wire _07048_;
 wire _07049_;
 wire _07050_;
 wire _07051_;
 wire _07052_;
 wire _07053_;
 wire _07054_;
 wire _07055_;
 wire _07056_;
 wire _07057_;
 wire _07058_;
 wire _07059_;
 wire _07060_;
 wire _07061_;
 wire _07062_;
 wire _07063_;
 wire _07064_;
 wire _07065_;
 wire _07066_;
 wire _07067_;
 wire _07068_;
 wire _07069_;
 wire _07070_;
 wire _07071_;
 wire _07072_;
 wire _07073_;
 wire _07074_;
 wire _07075_;
 wire _07076_;
 wire _07077_;
 wire _07078_;
 wire _07079_;
 wire _07080_;
 wire _07081_;
 wire _07082_;
 wire _07083_;
 wire _07084_;
 wire _07085_;
 wire _07086_;
 wire _07087_;
 wire _07088_;
 wire _07089_;
 wire _07090_;
 wire _07091_;
 wire _07092_;
 wire _07093_;
 wire _07094_;
 wire _07095_;
 wire _07096_;
 wire _07097_;
 wire _07098_;
 wire _07099_;
 wire _07100_;
 wire _07101_;
 wire _07102_;
 wire _07103_;
 wire _07104_;
 wire _07105_;
 wire _07106_;
 wire _07107_;
 wire _07108_;
 wire _07109_;
 wire _07110_;
 wire _07111_;
 wire _07112_;
 wire _07113_;
 wire _07114_;
 wire _07115_;
 wire _07116_;
 wire _07117_;
 wire _07118_;
 wire _07119_;
 wire _07120_;
 wire _07121_;
 wire _07122_;
 wire _07123_;
 wire _07124_;
 wire _07125_;
 wire _07126_;
 wire _07127_;
 wire _07128_;
 wire _07129_;
 wire _07130_;
 wire _07131_;
 wire _07132_;
 wire _07133_;
 wire _07134_;
 wire _07135_;
 wire _07136_;
 wire _07137_;
 wire _07138_;
 wire _07139_;
 wire _07140_;
 wire _07141_;
 wire _07142_;
 wire _07143_;
 wire _07144_;
 wire _07145_;
 wire _07146_;
 wire _07147_;
 wire _07148_;
 wire _07149_;
 wire _07150_;
 wire _07151_;
 wire _07152_;
 wire _07153_;
 wire _07154_;
 wire _07155_;
 wire _07156_;
 wire _07157_;
 wire _07158_;
 wire _07159_;
 wire _07160_;
 wire _07161_;
 wire _07162_;
 wire _07163_;
 wire _07164_;
 wire _07165_;
 wire _07166_;
 wire _07167_;
 wire _07168_;
 wire _07169_;
 wire _07170_;
 wire _07171_;
 wire _07172_;
 wire _07173_;
 wire _07174_;
 wire _07175_;
 wire _07176_;
 wire _07177_;
 wire _07178_;
 wire _07179_;
 wire _07180_;
 wire _07181_;
 wire _07182_;
 wire _07183_;
 wire _07184_;
 wire _07185_;
 wire _07186_;
 wire _07187_;
 wire _07188_;
 wire _07189_;
 wire _07190_;
 wire _07191_;
 wire _07192_;
 wire _07193_;
 wire _07194_;
 wire _07195_;
 wire _07196_;
 wire _07197_;
 wire _07198_;
 wire _07199_;
 wire _07200_;
 wire _07201_;
 wire _07202_;
 wire _07203_;
 wire _07204_;
 wire _07205_;
 wire _07206_;
 wire _07207_;
 wire _07208_;
 wire _07209_;
 wire _07210_;
 wire _07211_;
 wire _07212_;
 wire _07213_;
 wire _07214_;
 wire _07215_;
 wire _07216_;
 wire _07217_;
 wire _07218_;
 wire _07219_;
 wire _07220_;
 wire _07221_;
 wire _07222_;
 wire _07223_;
 wire _07224_;
 wire _07225_;
 wire _07226_;
 wire _07227_;
 wire _07228_;
 wire _07229_;
 wire _07230_;
 wire _07231_;
 wire _07232_;
 wire _07233_;
 wire _07234_;
 wire _07235_;
 wire _07236_;
 wire _07237_;
 wire _07238_;
 wire _07239_;
 wire _07240_;
 wire _07241_;
 wire _07242_;
 wire _07243_;
 wire _07244_;
 wire _07245_;
 wire _07246_;
 wire _07247_;
 wire _07248_;
 wire _07249_;
 wire _07250_;
 wire _07251_;
 wire _07252_;
 wire _07253_;
 wire _07254_;
 wire _07255_;
 wire _07256_;
 wire _07257_;
 wire _07258_;
 wire _07259_;
 wire _07260_;
 wire _07261_;
 wire _07262_;
 wire _07263_;
 wire _07264_;
 wire _07265_;
 wire _07266_;
 wire _07267_;
 wire _07268_;
 wire _07269_;
 wire _07270_;
 wire _07271_;
 wire _07272_;
 wire _07273_;
 wire _07274_;
 wire _07275_;
 wire _07276_;
 wire _07277_;
 wire _07278_;
 wire _07279_;
 wire _07280_;
 wire _07281_;
 wire _07282_;
 wire _07283_;
 wire _07284_;
 wire _07285_;
 wire _07286_;
 wire _07287_;
 wire _07288_;
 wire _07289_;
 wire _07290_;
 wire _07291_;
 wire _07292_;
 wire _07293_;
 wire _07294_;
 wire _07295_;
 wire _07296_;
 wire _07297_;
 wire _07298_;
 wire _07299_;
 wire _07300_;
 wire _07301_;
 wire _07302_;
 wire _07303_;
 wire _07304_;
 wire _07305_;
 wire _07306_;
 wire _07307_;
 wire _07308_;
 wire _07309_;
 wire _07310_;
 wire _07311_;
 wire _07312_;
 wire _07313_;
 wire _07314_;
 wire _07315_;
 wire _07316_;
 wire _07317_;
 wire _07318_;
 wire _07319_;
 wire _07320_;
 wire _07321_;
 wire _07322_;
 wire _07323_;
 wire _07324_;
 wire _07325_;
 wire _07326_;
 wire _07327_;
 wire _07328_;
 wire _07329_;
 wire _07330_;
 wire _07331_;
 wire _07332_;
 wire _07333_;
 wire _07334_;
 wire _07335_;
 wire _07336_;
 wire _07337_;
 wire _07338_;
 wire _07339_;
 wire _07340_;
 wire _07341_;
 wire _07342_;
 wire _07343_;
 wire _07344_;
 wire _07345_;
 wire _07346_;
 wire _07347_;
 wire _07348_;
 wire _07349_;
 wire _07350_;
 wire _07351_;
 wire _07352_;
 wire _07353_;
 wire _07354_;
 wire _07355_;
 wire _07356_;
 wire _07357_;
 wire _07358_;
 wire _07359_;
 wire _07360_;
 wire _07361_;
 wire _07362_;
 wire _07363_;
 wire _07364_;
 wire _07365_;
 wire _07366_;
 wire _07367_;
 wire _07368_;
 wire _07369_;
 wire _07370_;
 wire _07371_;
 wire _07372_;
 wire _07373_;
 wire _07374_;
 wire _07375_;
 wire _07376_;
 wire _07377_;
 wire _07378_;
 wire _07379_;
 wire _07380_;
 wire _07381_;
 wire _07382_;
 wire _07383_;
 wire _07384_;
 wire _07385_;
 wire _07386_;
 wire _07387_;
 wire _07388_;
 wire _07389_;
 wire _07390_;
 wire _07391_;
 wire _07392_;
 wire _07393_;
 wire _07394_;
 wire _07395_;
 wire _07396_;
 wire _07397_;
 wire _07398_;
 wire _07399_;
 wire _07400_;
 wire _07401_;
 wire _07402_;
 wire _07403_;
 wire _07404_;
 wire _07405_;
 wire net1239;
 wire _07407_;
 wire net66;
 wire _07409_;
 wire _07410_;
 wire _07411_;
 wire _07412_;
 wire _07413_;
 wire _07414_;
 wire _07415_;
 wire _07416_;
 wire _07417_;
 wire _07418_;
 wire _07419_;
 wire net18;
 wire _07421_;
 wire _07422_;
 wire _07423_;
 wire _07424_;
 wire _07425_;
 wire _07426_;
 wire _07427_;
 wire _07428_;
 wire _07429_;
 wire _07430_;
 wire _07431_;
 wire _07432_;
 wire _07433_;
 wire _07434_;
 wire _07435_;
 wire net28;
 wire _07437_;
 wire _07438_;
 wire _07439_;
 wire _07440_;
 wire _07441_;
 wire _07442_;
 wire _07443_;
 wire _07444_;
 wire _07445_;
 wire _07446_;
 wire _07447_;
 wire _07448_;
 wire _07449_;
 wire _07450_;
 wire _07451_;
 wire _07452_;
 wire _07453_;
 wire _07454_;
 wire _07455_;
 wire _07456_;
 wire _07457_;
 wire _07458_;
 wire _07459_;
 wire _07460_;
 wire _07461_;
 wire _07462_;
 wire _07463_;
 wire _07464_;
 wire _07465_;
 wire _07466_;
 wire _07467_;
 wire _07468_;
 wire _07469_;
 wire _07470_;
 wire net39;
 wire _07472_;
 wire _07473_;
 wire _07474_;
 wire _07475_;
 wire _07476_;
 wire _07477_;
 wire _07478_;
 wire _07479_;
 wire _07480_;
 wire _07481_;
 wire _07482_;
 wire _07483_;
 wire _07484_;
 wire _07485_;
 wire _07486_;
 wire _07487_;
 wire _07488_;
 wire _07489_;
 wire _07490_;
 wire _07491_;
 wire _07492_;
 wire _07493_;
 wire _07494_;
 wire _07495_;
 wire _07496_;
 wire _07497_;
 wire _07498_;
 wire _07499_;
 wire _07500_;
 wire _07501_;
 wire _07502_;
 wire _07503_;
 wire _07504_;
 wire _07505_;
 wire _07506_;
 wire _07507_;
 wire _07508_;
 wire _07509_;
 wire _07510_;
 wire _07511_;
 wire _07512_;
 wire _07513_;
 wire _07514_;
 wire _07515_;
 wire _07516_;
 wire _07517_;
 wire _07518_;
 wire _07519_;
 wire _07520_;
 wire _07521_;
 wire _07522_;
 wire _07523_;
 wire _07524_;
 wire _07525_;
 wire _07526_;
 wire _07527_;
 wire _07528_;
 wire _07529_;
 wire _07530_;
 wire _07531_;
 wire _07532_;
 wire _07533_;
 wire _07534_;
 wire _07535_;
 wire _07536_;
 wire _07537_;
 wire _07538_;
 wire _07539_;
 wire _07540_;
 wire _07541_;
 wire _07542_;
 wire _07543_;
 wire _07544_;
 wire _07545_;
 wire _07546_;
 wire _07547_;
 wire _07548_;
 wire _07549_;
 wire _07550_;
 wire _07551_;
 wire _07552_;
 wire _07553_;
 wire _07554_;
 wire _07555_;
 wire _07556_;
 wire _07557_;
 wire _07558_;
 wire _07559_;
 wire _07560_;
 wire _07561_;
 wire _07562_;
 wire _07563_;
 wire _07564_;
 wire _07565_;
 wire _07566_;
 wire _07567_;
 wire _07568_;
 wire _07569_;
 wire _07570_;
 wire _07571_;
 wire _07572_;
 wire _07573_;
 wire _07574_;
 wire _07575_;
 wire _07576_;
 wire _07577_;
 wire _07578_;
 wire _07579_;
 wire _07580_;
 wire _07581_;
 wire _07582_;
 wire _07583_;
 wire _07584_;
 wire _07585_;
 wire _07586_;
 wire _07587_;
 wire _07588_;
 wire _07589_;
 wire _07590_;
 wire _07591_;
 wire _07592_;
 wire _07593_;
 wire _07594_;
 wire _07595_;
 wire _07596_;
 wire _07597_;
 wire _07598_;
 wire _07599_;
 wire _07600_;
 wire _07601_;
 wire _07602_;
 wire _07603_;
 wire _07604_;
 wire _07605_;
 wire _07606_;
 wire _07607_;
 wire _07608_;
 wire _07609_;
 wire _07610_;
 wire _07611_;
 wire _07612_;
 wire _07613_;
 wire _07614_;
 wire _07615_;
 wire _07616_;
 wire _07617_;
 wire _07618_;
 wire _07619_;
 wire _07620_;
 wire _07621_;
 wire _07622_;
 wire _07623_;
 wire _07624_;
 wire _07625_;
 wire _07626_;
 wire _07627_;
 wire _07628_;
 wire _07629_;
 wire _07630_;
 wire _07631_;
 wire _07632_;
 wire _07633_;
 wire _07634_;
 wire _07635_;
 wire _07636_;
 wire _07637_;
 wire _07638_;
 wire _07639_;
 wire _07640_;
 wire _07641_;
 wire _07642_;
 wire _07643_;
 wire _07644_;
 wire _07645_;
 wire _07646_;
 wire _07647_;
 wire _07648_;
 wire _07649_;
 wire _07650_;
 wire _07651_;
 wire _07652_;
 wire _07653_;
 wire _07654_;
 wire _07655_;
 wire _07656_;
 wire _07657_;
 wire _07658_;
 wire _07659_;
 wire _07660_;
 wire _07661_;
 wire _07662_;
 wire _07663_;
 wire _07664_;
 wire _07665_;
 wire _07666_;
 wire _07667_;
 wire _07668_;
 wire _07669_;
 wire _07670_;
 wire _07671_;
 wire _07672_;
 wire _07673_;
 wire _07674_;
 wire _07675_;
 wire _07676_;
 wire _07677_;
 wire _07678_;
 wire _07679_;
 wire _07680_;
 wire _07681_;
 wire _07682_;
 wire _07683_;
 wire _07684_;
 wire _07685_;
 wire _07686_;
 wire _07687_;
 wire _07688_;
 wire _07689_;
 wire _07690_;
 wire _07691_;
 wire _07692_;
 wire _07693_;
 wire _07694_;
 wire _07695_;
 wire _07696_;
 wire _07697_;
 wire _07698_;
 wire _07699_;
 wire _07700_;
 wire _07701_;
 wire _07702_;
 wire _07703_;
 wire _07704_;
 wire _07705_;
 wire _07706_;
 wire _07707_;
 wire _07708_;
 wire _07709_;
 wire _07710_;
 wire _07711_;
 wire _07712_;
 wire _07713_;
 wire _07714_;
 wire _07715_;
 wire _07716_;
 wire _07717_;
 wire _07718_;
 wire _07719_;
 wire _07720_;
 wire _07721_;
 wire _07722_;
 wire _07723_;
 wire _07724_;
 wire _07725_;
 wire _07726_;
 wire _07727_;
 wire _07728_;
 wire _07729_;
 wire _07730_;
 wire _07731_;
 wire _07732_;
 wire _07733_;
 wire _07734_;
 wire _07735_;
 wire _07736_;
 wire _07737_;
 wire _07738_;
 wire _07739_;
 wire _07740_;
 wire _07741_;
 wire _07742_;
 wire _07743_;
 wire _07744_;
 wire _07745_;
 wire _07746_;
 wire _07747_;
 wire _07748_;
 wire _07749_;
 wire _07750_;
 wire _07751_;
 wire _07752_;
 wire _07753_;
 wire _07754_;
 wire _07755_;
 wire _07756_;
 wire _07757_;
 wire _07758_;
 wire _07759_;
 wire _07760_;
 wire _07761_;
 wire _07762_;
 wire _07763_;
 wire _07764_;
 wire _07765_;
 wire _07766_;
 wire _07767_;
 wire _07768_;
 wire _07769_;
 wire _07770_;
 wire _07771_;
 wire _07772_;
 wire _07773_;
 wire _07774_;
 wire _07775_;
 wire _07776_;
 wire _07777_;
 wire _07778_;
 wire _07779_;
 wire _07780_;
 wire _07781_;
 wire _07782_;
 wire _07783_;
 wire _07784_;
 wire _07785_;
 wire _07786_;
 wire _07787_;
 wire _07788_;
 wire _07789_;
 wire _07790_;
 wire _07791_;
 wire _07792_;
 wire _07793_;
 wire _07794_;
 wire _07795_;
 wire _07796_;
 wire _07797_;
 wire _07798_;
 wire _07799_;
 wire _07800_;
 wire _07801_;
 wire _07802_;
 wire _07803_;
 wire _07804_;
 wire _07805_;
 wire _07806_;
 wire _07807_;
 wire _07808_;
 wire _07809_;
 wire _07810_;
 wire _07811_;
 wire _07812_;
 wire _07813_;
 wire _07814_;
 wire _07815_;
 wire _07816_;
 wire _07817_;
 wire _07818_;
 wire _07819_;
 wire _07820_;
 wire _07821_;
 wire _07822_;
 wire _07823_;
 wire _07824_;
 wire _07825_;
 wire _07826_;
 wire _07827_;
 wire _07828_;
 wire _07829_;
 wire _07830_;
 wire _07831_;
 wire _07832_;
 wire _07833_;
 wire _07834_;
 wire _07835_;
 wire _07836_;
 wire _07837_;
 wire _07838_;
 wire _07839_;
 wire _07840_;
 wire _07841_;
 wire _07842_;
 wire _07843_;
 wire _07844_;
 wire _07845_;
 wire _07846_;
 wire _07847_;
 wire _07848_;
 wire _07849_;
 wire _07850_;
 wire _07851_;
 wire _07852_;
 wire _07853_;
 wire _07854_;
 wire _07855_;
 wire _07856_;
 wire _07857_;
 wire _07858_;
 wire _07859_;
 wire _07860_;
 wire _07861_;
 wire _07862_;
 wire _07863_;
 wire _07864_;
 wire _07865_;
 wire _07866_;
 wire _07867_;
 wire _07868_;
 wire _07869_;
 wire _07870_;
 wire _07871_;
 wire _07872_;
 wire _07873_;
 wire _07874_;
 wire _07875_;
 wire _07876_;
 wire _07877_;
 wire _07878_;
 wire _07879_;
 wire _07880_;
 wire _07881_;
 wire _07882_;
 wire _07883_;
 wire _07884_;
 wire _07885_;
 wire _07886_;
 wire _07887_;
 wire _07888_;
 wire _07889_;
 wire _07890_;
 wire _07891_;
 wire _07892_;
 wire _07893_;
 wire _07894_;
 wire _07895_;
 wire _07896_;
 wire _07897_;
 wire _07898_;
 wire _07899_;
 wire _07900_;
 wire _07901_;
 wire _07902_;
 wire _07903_;
 wire _07904_;
 wire _07905_;
 wire _07906_;
 wire _07907_;
 wire _07908_;
 wire _07909_;
 wire _07910_;
 wire _07911_;
 wire _07912_;
 wire _07913_;
 wire _07914_;
 wire _07915_;
 wire _07916_;
 wire _07917_;
 wire _07918_;
 wire _07919_;
 wire _07920_;
 wire _07921_;
 wire _07922_;
 wire _07923_;
 wire _07924_;
 wire _07925_;
 wire _07926_;
 wire _07927_;
 wire _07928_;
 wire _07929_;
 wire _07930_;
 wire _07931_;
 wire net101;
 wire _07933_;
 wire _07934_;
 wire _07935_;
 wire _07936_;
 wire _07937_;
 wire _07938_;
 wire _07939_;
 wire _07940_;
 wire _07941_;
 wire _07942_;
 wire _07943_;
 wire _07944_;
 wire net27;
 wire _07946_;
 wire _07947_;
 wire _07948_;
 wire _07949_;
 wire _07950_;
 wire net99;
 wire _07952_;
 wire _07953_;
 wire _07954_;
 wire _07955_;
 wire _07956_;
 wire _07957_;
 wire _07958_;
 wire _07959_;
 wire _07960_;
 wire _07961_;
 wire _07962_;
 wire _07963_;
 wire _07964_;
 wire _07965_;
 wire _07966_;
 wire _07967_;
 wire _07968_;
 wire _07969_;
 wire _07970_;
 wire _07971_;
 wire _07972_;
 wire _07973_;
 wire _07974_;
 wire _07975_;
 wire _07976_;
 wire _07977_;
 wire _07978_;
 wire _07979_;
 wire net1211;
 wire _07981_;
 wire _07982_;
 wire _07983_;
 wire _07984_;
 wire _07985_;
 wire _07986_;
 wire _07987_;
 wire _07988_;
 wire _07989_;
 wire _07990_;
 wire _07991_;
 wire _07992_;
 wire _07993_;
 wire _07994_;
 wire _07995_;
 wire _07996_;
 wire _07997_;
 wire _07998_;
 wire _07999_;
 wire _08000_;
 wire _08001_;
 wire _08002_;
 wire _08003_;
 wire _08004_;
 wire _08005_;
 wire _08006_;
 wire _08007_;
 wire _08008_;
 wire _08009_;
 wire _08010_;
 wire _08011_;
 wire _08012_;
 wire _08013_;
 wire _08014_;
 wire _08015_;
 wire _08016_;
 wire _08017_;
 wire _08018_;
 wire _08019_;
 wire _08020_;
 wire _08021_;
 wire _08022_;
 wire _08023_;
 wire _08024_;
 wire _08025_;
 wire _08026_;
 wire _08027_;
 wire _08028_;
 wire _08029_;
 wire _08030_;
 wire _08031_;
 wire _08032_;
 wire _08033_;
 wire _08034_;
 wire _08035_;
 wire _08036_;
 wire _08037_;
 wire _08038_;
 wire _08039_;
 wire _08040_;
 wire _08041_;
 wire _08042_;
 wire _08043_;
 wire _08044_;
 wire _08045_;
 wire _08046_;
 wire _08047_;
 wire _08048_;
 wire _08049_;
 wire _08050_;
 wire _08051_;
 wire _08052_;
 wire _08053_;
 wire _08054_;
 wire _08055_;
 wire _08056_;
 wire _08057_;
 wire _08058_;
 wire _08059_;
 wire _08060_;
 wire _08061_;
 wire _08062_;
 wire _08063_;
 wire _08064_;
 wire _08065_;
 wire _08066_;
 wire _08067_;
 wire _08068_;
 wire _08069_;
 wire _08070_;
 wire _08071_;
 wire _08072_;
 wire _08073_;
 wire _08074_;
 wire _08075_;
 wire _08076_;
 wire _08077_;
 wire _08078_;
 wire _08079_;
 wire _08080_;
 wire _08081_;
 wire _08082_;
 wire _08083_;
 wire _08084_;
 wire _08085_;
 wire _08086_;
 wire _08087_;
 wire _08088_;
 wire _08089_;
 wire _08090_;
 wire _08091_;
 wire _08092_;
 wire _08093_;
 wire _08094_;
 wire _08095_;
 wire _08096_;
 wire _08097_;
 wire _08098_;
 wire _08099_;
 wire _08100_;
 wire _08101_;
 wire _08102_;
 wire _08103_;
 wire _08104_;
 wire _08105_;
 wire _08106_;
 wire _08107_;
 wire _08108_;
 wire _08109_;
 wire _08110_;
 wire _08111_;
 wire _08112_;
 wire _08113_;
 wire _08114_;
 wire _08115_;
 wire _08116_;
 wire _08117_;
 wire _08118_;
 wire _08119_;
 wire _08120_;
 wire _08121_;
 wire _08122_;
 wire _08123_;
 wire _08124_;
 wire _08125_;
 wire _08126_;
 wire _08127_;
 wire _08128_;
 wire _08129_;
 wire _08130_;
 wire _08131_;
 wire _08132_;
 wire _08133_;
 wire _08134_;
 wire _08135_;
 wire _08136_;
 wire _08137_;
 wire _08138_;
 wire _08139_;
 wire _08140_;
 wire _08141_;
 wire _08142_;
 wire _08143_;
 wire _08144_;
 wire _08145_;
 wire _08146_;
 wire _08147_;
 wire _08148_;
 wire _08149_;
 wire _08150_;
 wire _08151_;
 wire _08152_;
 wire _08153_;
 wire _08154_;
 wire _08155_;
 wire _08156_;
 wire _08157_;
 wire _08158_;
 wire _08159_;
 wire _08160_;
 wire _08161_;
 wire _08162_;
 wire _08163_;
 wire _08164_;
 wire _08165_;
 wire _08166_;
 wire _08167_;
 wire _08168_;
 wire _08169_;
 wire _08170_;
 wire _08171_;
 wire _08172_;
 wire _08173_;
 wire _08174_;
 wire _08175_;
 wire _08176_;
 wire _08177_;
 wire _08178_;
 wire _08179_;
 wire _08180_;
 wire _08181_;
 wire _08182_;
 wire _08183_;
 wire _08184_;
 wire _08185_;
 wire _08186_;
 wire _08187_;
 wire _08188_;
 wire _08189_;
 wire _08190_;
 wire _08191_;
 wire _08192_;
 wire _08193_;
 wire _08194_;
 wire _08195_;
 wire _08196_;
 wire _08197_;
 wire _08198_;
 wire _08199_;
 wire _08200_;
 wire _08201_;
 wire _08202_;
 wire _08203_;
 wire _08204_;
 wire _08205_;
 wire _08206_;
 wire _08207_;
 wire _08208_;
 wire _08209_;
 wire _08210_;
 wire _08211_;
 wire _08212_;
 wire _08213_;
 wire _08214_;
 wire _08215_;
 wire _08216_;
 wire _08217_;
 wire _08218_;
 wire _08219_;
 wire _08220_;
 wire _08221_;
 wire _08222_;
 wire _08223_;
 wire _08224_;
 wire _08225_;
 wire _08226_;
 wire _08227_;
 wire _08228_;
 wire _08229_;
 wire _08230_;
 wire _08231_;
 wire _08232_;
 wire _08233_;
 wire _08234_;
 wire _08235_;
 wire _08236_;
 wire _08237_;
 wire _08238_;
 wire _08239_;
 wire _08240_;
 wire _08241_;
 wire _08242_;
 wire _08243_;
 wire _08244_;
 wire _08245_;
 wire _08246_;
 wire _08247_;
 wire _08248_;
 wire _08249_;
 wire _08250_;
 wire _08251_;
 wire _08252_;
 wire _08253_;
 wire _08254_;
 wire _08255_;
 wire _08256_;
 wire _08257_;
 wire _08258_;
 wire _08259_;
 wire _08260_;
 wire _08261_;
 wire _08262_;
 wire _08263_;
 wire _08264_;
 wire _08265_;
 wire _08266_;
 wire _08267_;
 wire _08268_;
 wire _08269_;
 wire _08270_;
 wire _08271_;
 wire _08272_;
 wire _08273_;
 wire _08274_;
 wire _08275_;
 wire _08276_;
 wire _08277_;
 wire _08278_;
 wire _08279_;
 wire _08280_;
 wire _08281_;
 wire _08282_;
 wire _08283_;
 wire _08284_;
 wire _08285_;
 wire _08286_;
 wire _08287_;
 wire _08288_;
 wire _08289_;
 wire _08290_;
 wire _08291_;
 wire _08292_;
 wire _08293_;
 wire _08294_;
 wire _08295_;
 wire _08296_;
 wire _08297_;
 wire _08298_;
 wire _08299_;
 wire _08300_;
 wire _08301_;
 wire _08302_;
 wire _08303_;
 wire _08304_;
 wire _08305_;
 wire _08306_;
 wire _08307_;
 wire _08308_;
 wire _08309_;
 wire _08310_;
 wire _08311_;
 wire _08312_;
 wire _08313_;
 wire _08314_;
 wire _08315_;
 wire _08316_;
 wire _08317_;
 wire _08318_;
 wire _08319_;
 wire _08320_;
 wire _08321_;
 wire _08322_;
 wire _08323_;
 wire _08324_;
 wire _08325_;
 wire _08326_;
 wire _08327_;
 wire _08328_;
 wire _08329_;
 wire _08330_;
 wire _08331_;
 wire _08332_;
 wire _08333_;
 wire _08334_;
 wire _08335_;
 wire _08336_;
 wire _08337_;
 wire _08338_;
 wire _08339_;
 wire _08340_;
 wire _08341_;
 wire _08342_;
 wire _08343_;
 wire _08344_;
 wire _08345_;
 wire _08346_;
 wire _08347_;
 wire _08348_;
 wire _08349_;
 wire _08350_;
 wire _08351_;
 wire _08352_;
 wire _08353_;
 wire _08354_;
 wire _08355_;
 wire _08356_;
 wire _08357_;
 wire _08358_;
 wire _08359_;
 wire _08360_;
 wire _08361_;
 wire _08362_;
 wire _08363_;
 wire _08364_;
 wire _08365_;
 wire _08366_;
 wire _08367_;
 wire _08368_;
 wire _08369_;
 wire _08370_;
 wire _08371_;
 wire _08372_;
 wire _08373_;
 wire _08374_;
 wire _08375_;
 wire _08376_;
 wire _08377_;
 wire _08378_;
 wire _08379_;
 wire _08380_;
 wire _08381_;
 wire _08382_;
 wire _08383_;
 wire _08384_;
 wire _08385_;
 wire _08386_;
 wire _08387_;
 wire _08388_;
 wire _08389_;
 wire _08390_;
 wire _08391_;
 wire _08392_;
 wire _08393_;
 wire _08394_;
 wire _08395_;
 wire _08396_;
 wire _08397_;
 wire _08398_;
 wire _08399_;
 wire _08400_;
 wire _08401_;
 wire _08402_;
 wire _08403_;
 wire _08404_;
 wire _08405_;
 wire _08406_;
 wire _08407_;
 wire _08408_;
 wire _08409_;
 wire _08410_;
 wire _08411_;
 wire _08412_;
 wire _08413_;
 wire _08414_;
 wire _08415_;
 wire _08416_;
 wire _08417_;
 wire _08418_;
 wire _08419_;
 wire _08420_;
 wire _08421_;
 wire _08422_;
 wire _08423_;
 wire _08424_;
 wire _08425_;
 wire _08426_;
 wire _08427_;
 wire _08428_;
 wire _08429_;
 wire _08430_;
 wire _08431_;
 wire _08432_;
 wire _08433_;
 wire _08434_;
 wire _08435_;
 wire _08436_;
 wire _08437_;
 wire _08438_;
 wire _08439_;
 wire _08440_;
 wire _08441_;
 wire _08442_;
 wire _08443_;
 wire net51;
 wire _08445_;
 wire _08446_;
 wire _08447_;
 wire _08448_;
 wire _08449_;
 wire _08450_;
 wire net1127;
 wire _08452_;
 wire _08453_;
 wire _08454_;
 wire _08455_;
 wire _08456_;
 wire _08457_;
 wire _08458_;
 wire _08459_;
 wire _08460_;
 wire _08461_;
 wire _08462_;
 wire _08463_;
 wire _08464_;
 wire _08465_;
 wire _08466_;
 wire _08467_;
 wire _08468_;
 wire _08469_;
 wire _08470_;
 wire _08471_;
 wire _08472_;
 wire _08473_;
 wire _08474_;
 wire _08475_;
 wire net100;
 wire _08477_;
 wire _08478_;
 wire _08479_;
 wire _08480_;
 wire _08481_;
 wire _08482_;
 wire _08483_;
 wire _08484_;
 wire _08485_;
 wire _08486_;
 wire _08487_;
 wire _08488_;
 wire _08489_;
 wire _08490_;
 wire _08491_;
 wire _08492_;
 wire _08493_;
 wire _08494_;
 wire _08495_;
 wire _08496_;
 wire _08497_;
 wire _08498_;
 wire _08499_;
 wire _08500_;
 wire _08501_;
 wire _08502_;
 wire _08503_;
 wire _08504_;
 wire _08505_;
 wire _08506_;
 wire _08507_;
 wire _08508_;
 wire _08509_;
 wire _08510_;
 wire _08511_;
 wire _08512_;
 wire _08513_;
 wire _08514_;
 wire _08515_;
 wire _08516_;
 wire _08517_;
 wire _08518_;
 wire _08519_;
 wire _08520_;
 wire _08521_;
 wire _08522_;
 wire _08523_;
 wire _08524_;
 wire _08525_;
 wire _08526_;
 wire _08527_;
 wire _08528_;
 wire _08529_;
 wire _08530_;
 wire _08531_;
 wire _08532_;
 wire _08533_;
 wire _08534_;
 wire _08535_;
 wire _08536_;
 wire _08537_;
 wire _08538_;
 wire _08539_;
 wire _08540_;
 wire _08541_;
 wire _08542_;
 wire _08543_;
 wire _08544_;
 wire _08545_;
 wire _08546_;
 wire _08547_;
 wire _08548_;
 wire _08549_;
 wire _08550_;
 wire _08551_;
 wire _08552_;
 wire _08553_;
 wire _08554_;
 wire _08555_;
 wire _08556_;
 wire _08557_;
 wire _08558_;
 wire _08559_;
 wire _08560_;
 wire _08561_;
 wire _08562_;
 wire _08563_;
 wire _08564_;
 wire _08565_;
 wire _08566_;
 wire _08567_;
 wire _08568_;
 wire _08569_;
 wire _08570_;
 wire _08571_;
 wire _08572_;
 wire _08573_;
 wire _08574_;
 wire _08575_;
 wire _08576_;
 wire _08577_;
 wire _08578_;
 wire _08579_;
 wire _08580_;
 wire _08581_;
 wire _08582_;
 wire _08583_;
 wire _08584_;
 wire _08585_;
 wire _08586_;
 wire _08587_;
 wire _08588_;
 wire _08589_;
 wire _08590_;
 wire _08591_;
 wire _08592_;
 wire _08593_;
 wire _08594_;
 wire _08595_;
 wire _08596_;
 wire _08597_;
 wire _08598_;
 wire _08599_;
 wire _08600_;
 wire _08601_;
 wire _08602_;
 wire _08603_;
 wire _08604_;
 wire _08605_;
 wire _08606_;
 wire _08607_;
 wire _08608_;
 wire _08609_;
 wire _08610_;
 wire _08611_;
 wire _08612_;
 wire _08613_;
 wire _08614_;
 wire _08615_;
 wire _08616_;
 wire _08617_;
 wire _08618_;
 wire _08619_;
 wire _08620_;
 wire _08621_;
 wire _08622_;
 wire _08623_;
 wire _08624_;
 wire _08625_;
 wire _08626_;
 wire _08627_;
 wire _08628_;
 wire _08629_;
 wire _08630_;
 wire _08631_;
 wire _08632_;
 wire _08633_;
 wire _08634_;
 wire _08635_;
 wire _08636_;
 wire _08637_;
 wire _08638_;
 wire _08639_;
 wire _08640_;
 wire _08641_;
 wire _08642_;
 wire _08643_;
 wire _08644_;
 wire _08645_;
 wire _08646_;
 wire _08647_;
 wire _08648_;
 wire _08649_;
 wire _08650_;
 wire _08651_;
 wire _08652_;
 wire _08653_;
 wire _08654_;
 wire _08655_;
 wire _08656_;
 wire _08657_;
 wire _08658_;
 wire _08659_;
 wire _08660_;
 wire _08661_;
 wire _08662_;
 wire _08663_;
 wire _08664_;
 wire _08665_;
 wire _08666_;
 wire _08667_;
 wire _08668_;
 wire _08669_;
 wire _08670_;
 wire _08671_;
 wire _08672_;
 wire _08673_;
 wire _08674_;
 wire _08675_;
 wire _08676_;
 wire _08677_;
 wire _08678_;
 wire _08679_;
 wire _08680_;
 wire _08681_;
 wire _08682_;
 wire _08683_;
 wire _08684_;
 wire _08685_;
 wire _08686_;
 wire _08687_;
 wire _08688_;
 wire _08689_;
 wire _08690_;
 wire _08691_;
 wire _08692_;
 wire _08693_;
 wire _08694_;
 wire _08695_;
 wire _08696_;
 wire _08697_;
 wire _08698_;
 wire _08699_;
 wire _08700_;
 wire _08701_;
 wire _08702_;
 wire _08703_;
 wire _08704_;
 wire _08705_;
 wire _08706_;
 wire _08707_;
 wire _08708_;
 wire _08709_;
 wire _08710_;
 wire _08711_;
 wire _08712_;
 wire _08713_;
 wire _08714_;
 wire _08715_;
 wire _08716_;
 wire _08717_;
 wire _08718_;
 wire _08719_;
 wire _08720_;
 wire _08721_;
 wire _08722_;
 wire _08723_;
 wire _08724_;
 wire _08725_;
 wire _08726_;
 wire _08727_;
 wire _08728_;
 wire _08729_;
 wire _08730_;
 wire _08731_;
 wire _08732_;
 wire _08733_;
 wire _08734_;
 wire _08735_;
 wire _08736_;
 wire _08737_;
 wire _08738_;
 wire _08739_;
 wire _08740_;
 wire _08741_;
 wire _08742_;
 wire _08743_;
 wire _08744_;
 wire _08745_;
 wire _08746_;
 wire _08747_;
 wire _08748_;
 wire _08749_;
 wire _08750_;
 wire _08751_;
 wire _08752_;
 wire _08753_;
 wire _08754_;
 wire _08755_;
 wire _08756_;
 wire _08757_;
 wire _08758_;
 wire _08759_;
 wire _08760_;
 wire _08761_;
 wire _08762_;
 wire _08763_;
 wire _08764_;
 wire _08765_;
 wire _08766_;
 wire _08767_;
 wire _08768_;
 wire _08769_;
 wire _08770_;
 wire _08771_;
 wire _08772_;
 wire _08773_;
 wire _08774_;
 wire _08775_;
 wire _08776_;
 wire _08777_;
 wire _08778_;
 wire _08779_;
 wire _08780_;
 wire _08781_;
 wire _08782_;
 wire _08783_;
 wire _08784_;
 wire _08785_;
 wire _08786_;
 wire _08787_;
 wire _08788_;
 wire _08789_;
 wire _08790_;
 wire _08791_;
 wire _08792_;
 wire _08793_;
 wire _08794_;
 wire _08795_;
 wire _08796_;
 wire _08797_;
 wire _08798_;
 wire _08799_;
 wire _08800_;
 wire _08801_;
 wire _08802_;
 wire _08803_;
 wire _08804_;
 wire _08805_;
 wire _08806_;
 wire _08807_;
 wire _08808_;
 wire _08809_;
 wire _08810_;
 wire _08811_;
 wire _08812_;
 wire _08813_;
 wire _08814_;
 wire _08815_;
 wire _08816_;
 wire _08817_;
 wire _08818_;
 wire _08819_;
 wire _08820_;
 wire _08821_;
 wire _08822_;
 wire _08823_;
 wire _08824_;
 wire _08825_;
 wire _08826_;
 wire _08827_;
 wire _08828_;
 wire _08829_;
 wire _08830_;
 wire _08831_;
 wire _08832_;
 wire _08833_;
 wire _08834_;
 wire _08835_;
 wire _08836_;
 wire _08837_;
 wire _08838_;
 wire _08839_;
 wire _08840_;
 wire _08841_;
 wire _08842_;
 wire _08843_;
 wire _08844_;
 wire _08845_;
 wire _08846_;
 wire _08847_;
 wire _08848_;
 wire _08849_;
 wire _08850_;
 wire _08851_;
 wire _08852_;
 wire _08853_;
 wire _08854_;
 wire _08855_;
 wire _08856_;
 wire _08857_;
 wire _08858_;
 wire _08859_;
 wire _08860_;
 wire _08861_;
 wire _08862_;
 wire _08863_;
 wire _08864_;
 wire _08865_;
 wire _08866_;
 wire _08867_;
 wire _08868_;
 wire _08869_;
 wire _08870_;
 wire _08871_;
 wire _08872_;
 wire _08873_;
 wire _08874_;
 wire _08875_;
 wire _08876_;
 wire _08877_;
 wire _08878_;
 wire _08879_;
 wire _08880_;
 wire _08881_;
 wire _08882_;
 wire _08883_;
 wire _08884_;
 wire _08885_;
 wire _08886_;
 wire _08887_;
 wire _08888_;
 wire _08889_;
 wire _08890_;
 wire _08891_;
 wire _08892_;
 wire _08893_;
 wire _08894_;
 wire _08895_;
 wire _08896_;
 wire _08897_;
 wire _08898_;
 wire _08899_;
 wire _08900_;
 wire _08901_;
 wire _08902_;
 wire _08903_;
 wire _08904_;
 wire _08905_;
 wire _08906_;
 wire _08907_;
 wire _08908_;
 wire _08909_;
 wire _08910_;
 wire _08911_;
 wire _08912_;
 wire _08913_;
 wire _08914_;
 wire _08915_;
 wire _08916_;
 wire _08917_;
 wire _08918_;
 wire _08919_;
 wire _08920_;
 wire _08921_;
 wire _08922_;
 wire _08923_;
 wire _08924_;
 wire _08925_;
 wire _08926_;
 wire _08927_;
 wire _08928_;
 wire _08929_;
 wire _08930_;
 wire _08931_;
 wire _08932_;
 wire _08933_;
 wire _08934_;
 wire _08935_;
 wire _08936_;
 wire _08937_;
 wire _08938_;
 wire _08939_;
 wire _08940_;
 wire _08941_;
 wire _08942_;
 wire _08943_;
 wire _08944_;
 wire _08945_;
 wire _08946_;
 wire _08947_;
 wire _08948_;
 wire _08949_;
 wire _08950_;
 wire _08951_;
 wire _08952_;
 wire _08953_;
 wire _08954_;
 wire _08955_;
 wire _08956_;
 wire _08957_;
 wire _08958_;
 wire _08959_;
 wire _08960_;
 wire _08961_;
 wire _08962_;
 wire _08963_;
 wire _08964_;
 wire _08965_;
 wire _08966_;
 wire _08967_;
 wire _08968_;
 wire _08969_;
 wire _08970_;
 wire _08971_;
 wire _08972_;
 wire _08973_;
 wire _08974_;
 wire _08975_;
 wire _08976_;
 wire _08977_;
 wire _08978_;
 wire _08979_;
 wire _08980_;
 wire net29;
 wire net8;
 wire _08983_;
 wire _08984_;
 wire net36;
 wire _08986_;
 wire _08987_;
 wire _08988_;
 wire _08989_;
 wire _08990_;
 wire _08991_;
 wire _08992_;
 wire _08993_;
 wire _08994_;
 wire _08995_;
 wire _08996_;
 wire _08997_;
 wire _08998_;
 wire _08999_;
 wire _09000_;
 wire _09001_;
 wire _09002_;
 wire _09003_;
 wire net884;
 wire net37;
 wire _09006_;
 wire _09007_;
 wire _09008_;
 wire _09009_;
 wire _09010_;
 wire _09011_;
 wire _09012_;
 wire _09013_;
 wire _09014_;
 wire _09015_;
 wire _09016_;
 wire _09017_;
 wire _09018_;
 wire _09019_;
 wire _09020_;
 wire _09021_;
 wire _09022_;
 wire _09023_;
 wire _09024_;
 wire _09025_;
 wire _09026_;
 wire _09027_;
 wire _09028_;
 wire _09029_;
 wire _09030_;
 wire _09031_;
 wire _09032_;
 wire _09033_;
 wire _09034_;
 wire net1160;
 wire net16;
 wire _09037_;
 wire _09038_;
 wire _09039_;
 wire _09040_;
 wire _09041_;
 wire _09042_;
 wire _09043_;
 wire _09044_;
 wire _09045_;
 wire _09046_;
 wire _09047_;
 wire _09048_;
 wire _09049_;
 wire _09050_;
 wire _09051_;
 wire _09052_;
 wire _09053_;
 wire _09054_;
 wire _09055_;
 wire _09056_;
 wire _09057_;
 wire _09058_;
 wire _09059_;
 wire _09060_;
 wire _09061_;
 wire _09062_;
 wire _09063_;
 wire _09064_;
 wire _09065_;
 wire _09066_;
 wire _09067_;
 wire _09068_;
 wire _09069_;
 wire _09070_;
 wire _09071_;
 wire _09072_;
 wire _09073_;
 wire _09074_;
 wire _09075_;
 wire _09076_;
 wire _09077_;
 wire _09078_;
 wire _09079_;
 wire _09080_;
 wire _09081_;
 wire _09082_;
 wire _09083_;
 wire _09084_;
 wire _09085_;
 wire _09086_;
 wire _09087_;
 wire _09088_;
 wire _09089_;
 wire _09090_;
 wire _09091_;
 wire _09092_;
 wire _09093_;
 wire _09094_;
 wire _09095_;
 wire _09096_;
 wire _09097_;
 wire _09098_;
 wire _09099_;
 wire _09100_;
 wire _09101_;
 wire _09102_;
 wire _09103_;
 wire _09104_;
 wire _09105_;
 wire _09106_;
 wire _09107_;
 wire _09108_;
 wire _09109_;
 wire _09110_;
 wire _09111_;
 wire _09112_;
 wire _09113_;
 wire _09114_;
 wire _09115_;
 wire _09116_;
 wire _09117_;
 wire _09118_;
 wire _09119_;
 wire _09120_;
 wire _09121_;
 wire _09122_;
 wire _09123_;
 wire _09124_;
 wire _09125_;
 wire _09126_;
 wire _09127_;
 wire _09128_;
 wire _09129_;
 wire _09130_;
 wire _09131_;
 wire _09132_;
 wire _09133_;
 wire _09134_;
 wire _09135_;
 wire _09136_;
 wire _09137_;
 wire _09138_;
 wire _09139_;
 wire _09140_;
 wire _09141_;
 wire _09142_;
 wire _09143_;
 wire net122;
 wire _09145_;
 wire _09146_;
 wire _09147_;
 wire _09148_;
 wire _09149_;
 wire _09150_;
 wire _09151_;
 wire _09152_;
 wire _09153_;
 wire _09154_;
 wire _09155_;
 wire _09156_;
 wire _09157_;
 wire _09158_;
 wire _09159_;
 wire _09160_;
 wire _09161_;
 wire _09162_;
 wire _09163_;
 wire _09164_;
 wire _09165_;
 wire _09166_;
 wire _09167_;
 wire _09168_;
 wire _09169_;
 wire _09170_;
 wire _09171_;
 wire _09172_;
 wire _09173_;
 wire _09174_;
 wire _09175_;
 wire _09176_;
 wire _09177_;
 wire _09178_;
 wire _09179_;
 wire _09180_;
 wire _09181_;
 wire _09182_;
 wire _09183_;
 wire _09184_;
 wire _09185_;
 wire _09186_;
 wire _09187_;
 wire _09188_;
 wire _09189_;
 wire _09190_;
 wire _09191_;
 wire _09192_;
 wire _09193_;
 wire _09194_;
 wire _09195_;
 wire _09196_;
 wire _09197_;
 wire _09198_;
 wire _09199_;
 wire _09200_;
 wire _09201_;
 wire _09202_;
 wire _09203_;
 wire _09204_;
 wire _09205_;
 wire _09206_;
 wire _09207_;
 wire _09208_;
 wire _09209_;
 wire _09210_;
 wire _09211_;
 wire _09212_;
 wire _09213_;
 wire _09214_;
 wire _09215_;
 wire _09216_;
 wire _09217_;
 wire _09218_;
 wire _09219_;
 wire _09220_;
 wire _09221_;
 wire _09222_;
 wire _09223_;
 wire _09224_;
 wire _09225_;
 wire _09226_;
 wire _09227_;
 wire _09228_;
 wire _09229_;
 wire _09230_;
 wire _09231_;
 wire _09232_;
 wire _09233_;
 wire _09234_;
 wire _09235_;
 wire _09236_;
 wire _09237_;
 wire _09238_;
 wire _09239_;
 wire _09240_;
 wire _09241_;
 wire _09242_;
 wire _09243_;
 wire _09244_;
 wire _09245_;
 wire _09246_;
 wire _09247_;
 wire _09248_;
 wire _09249_;
 wire _09250_;
 wire _09251_;
 wire _09252_;
 wire _09253_;
 wire _09254_;
 wire _09255_;
 wire _09256_;
 wire _09257_;
 wire _09258_;
 wire _09259_;
 wire _09260_;
 wire _09261_;
 wire _09262_;
 wire _09263_;
 wire _09264_;
 wire _09265_;
 wire _09266_;
 wire _09267_;
 wire _09268_;
 wire _09269_;
 wire _09270_;
 wire _09271_;
 wire _09272_;
 wire _09273_;
 wire _09274_;
 wire _09275_;
 wire _09276_;
 wire _09277_;
 wire _09278_;
 wire _09279_;
 wire _09280_;
 wire _09281_;
 wire _09282_;
 wire _09283_;
 wire _09284_;
 wire _09285_;
 wire _09286_;
 wire _09287_;
 wire _09288_;
 wire _09289_;
 wire net662;
 wire _09291_;
 wire _09292_;
 wire _09293_;
 wire _09294_;
 wire _09295_;
 wire net93;
 wire _09297_;
 wire _09298_;
 wire _09299_;
 wire _09300_;
 wire _09301_;
 wire _09302_;
 wire _09303_;
 wire _09304_;
 wire _09305_;
 wire _09306_;
 wire _09307_;
 wire _09308_;
 wire _09309_;
 wire _09310_;
 wire _09311_;
 wire _09312_;
 wire _09313_;
 wire _09314_;
 wire _09315_;
 wire _09316_;
 wire _09317_;
 wire _09318_;
 wire _09319_;
 wire _09320_;
 wire _09321_;
 wire _09322_;
 wire _09323_;
 wire _09324_;
 wire _09325_;
 wire _09326_;
 wire _09327_;
 wire _09328_;
 wire _09329_;
 wire _09330_;
 wire _09331_;
 wire _09332_;
 wire _09333_;
 wire _09334_;
 wire _09335_;
 wire _09336_;
 wire _09337_;
 wire _09338_;
 wire _09339_;
 wire _09340_;
 wire _09341_;
 wire _09342_;
 wire _09343_;
 wire _09344_;
 wire _09345_;
 wire _09346_;
 wire _09347_;
 wire _09348_;
 wire _09349_;
 wire _09350_;
 wire _09351_;
 wire _09352_;
 wire _09353_;
 wire _09354_;
 wire _09355_;
 wire _09356_;
 wire _09357_;
 wire _09358_;
 wire _09359_;
 wire _09360_;
 wire _09361_;
 wire _09362_;
 wire _09363_;
 wire _09364_;
 wire _09365_;
 wire _09366_;
 wire _09367_;
 wire _09368_;
 wire _09369_;
 wire _09370_;
 wire _09371_;
 wire _09372_;
 wire _09373_;
 wire _09374_;
 wire _09375_;
 wire _09376_;
 wire _09377_;
 wire _09378_;
 wire _09379_;
 wire _09380_;
 wire _09381_;
 wire _09382_;
 wire _09383_;
 wire _09384_;
 wire _09385_;
 wire _09386_;
 wire _09387_;
 wire _09388_;
 wire _09389_;
 wire _09390_;
 wire _09391_;
 wire _09392_;
 wire _09393_;
 wire _09394_;
 wire _09395_;
 wire _09396_;
 wire _09397_;
 wire _09398_;
 wire _09399_;
 wire _09400_;
 wire _09401_;
 wire _09402_;
 wire _09403_;
 wire _09404_;
 wire _09405_;
 wire _09406_;
 wire _09407_;
 wire _09408_;
 wire _09409_;
 wire _09410_;
 wire _09411_;
 wire _09412_;
 wire _09413_;
 wire _09414_;
 wire _09415_;
 wire _09416_;
 wire _09417_;
 wire _09418_;
 wire _09419_;
 wire _09420_;
 wire _09421_;
 wire _09422_;
 wire _09423_;
 wire _09424_;
 wire _09425_;
 wire _09426_;
 wire _09427_;
 wire _09428_;
 wire _09429_;
 wire _09430_;
 wire _09431_;
 wire _09432_;
 wire _09433_;
 wire _09434_;
 wire _09435_;
 wire _09436_;
 wire _09437_;
 wire _09438_;
 wire _09439_;
 wire _09440_;
 wire _09441_;
 wire _09442_;
 wire _09443_;
 wire _09444_;
 wire _09445_;
 wire _09446_;
 wire _09447_;
 wire _09448_;
 wire _09449_;
 wire _09450_;
 wire _09451_;
 wire _09452_;
 wire _09453_;
 wire _09454_;
 wire _09455_;
 wire _09456_;
 wire _09457_;
 wire _09458_;
 wire _09459_;
 wire _09460_;
 wire _09461_;
 wire _09462_;
 wire _09463_;
 wire _09464_;
 wire _09465_;
 wire _09466_;
 wire _09467_;
 wire _09468_;
 wire _09469_;
 wire _09470_;
 wire _09471_;
 wire _09472_;
 wire _09473_;
 wire _09474_;
 wire _09475_;
 wire _09476_;
 wire _09477_;
 wire _09478_;
 wire _09479_;
 wire _09480_;
 wire _09481_;
 wire _09482_;
 wire _09483_;
 wire _09484_;
 wire _09485_;
 wire _09486_;
 wire _09487_;
 wire _09488_;
 wire _09489_;
 wire _09490_;
 wire _09491_;
 wire _09492_;
 wire _09493_;
 wire _09494_;
 wire _09495_;
 wire _09496_;
 wire _09497_;
 wire _09498_;
 wire _09499_;
 wire _09500_;
 wire _09501_;
 wire _09502_;
 wire _09503_;
 wire _09504_;
 wire _09505_;
 wire _09506_;
 wire _09507_;
 wire _09508_;
 wire _09509_;
 wire _09510_;
 wire _09511_;
 wire _09512_;
 wire _09513_;
 wire _09514_;
 wire _09515_;
 wire _09516_;
 wire _09517_;
 wire _09518_;
 wire _09519_;
 wire _09520_;
 wire _09521_;
 wire _09522_;
 wire _09523_;
 wire _09524_;
 wire _09525_;
 wire _09526_;
 wire _09527_;
 wire _09528_;
 wire _09529_;
 wire _09530_;
 wire _09531_;
 wire _09532_;
 wire _09533_;
 wire _09534_;
 wire _09535_;
 wire _09536_;
 wire _09537_;
 wire _09538_;
 wire _09539_;
 wire _09540_;
 wire _09541_;
 wire _09542_;
 wire _09543_;
 wire _09544_;
 wire _09545_;
 wire _09546_;
 wire _09547_;
 wire _09548_;
 wire _09549_;
 wire _09550_;
 wire _09551_;
 wire _09552_;
 wire _09553_;
 wire _09554_;
 wire _09555_;
 wire _09556_;
 wire _09557_;
 wire _09558_;
 wire _09559_;
 wire _09560_;
 wire _09561_;
 wire _09562_;
 wire _09563_;
 wire _09564_;
 wire _09565_;
 wire _09566_;
 wire _09567_;
 wire _09568_;
 wire _09569_;
 wire _09570_;
 wire _09571_;
 wire _09572_;
 wire _09573_;
 wire _09574_;
 wire _09575_;
 wire _09576_;
 wire _09577_;
 wire _09578_;
 wire _09579_;
 wire _09580_;
 wire _09581_;
 wire _09582_;
 wire _09583_;
 wire _09584_;
 wire _09585_;
 wire _09586_;
 wire _09587_;
 wire _09588_;
 wire _09589_;
 wire _09590_;
 wire _09591_;
 wire _09592_;
 wire _09593_;
 wire _09594_;
 wire _09595_;
 wire _09596_;
 wire _09597_;
 wire _09598_;
 wire _09599_;
 wire _09600_;
 wire _09601_;
 wire _09602_;
 wire _09603_;
 wire _09604_;
 wire _09605_;
 wire _09606_;
 wire _09607_;
 wire _09608_;
 wire _09609_;
 wire _09610_;
 wire _09611_;
 wire _09612_;
 wire _09613_;
 wire _09614_;
 wire _09615_;
 wire _09616_;
 wire _09617_;
 wire _09618_;
 wire _09619_;
 wire _09620_;
 wire _09621_;
 wire _09622_;
 wire _09623_;
 wire _09624_;
 wire _09625_;
 wire _09626_;
 wire _09627_;
 wire _09628_;
 wire _09629_;
 wire _09630_;
 wire _09631_;
 wire _09632_;
 wire _09633_;
 wire _09634_;
 wire _09635_;
 wire _09636_;
 wire _09637_;
 wire _09638_;
 wire _09639_;
 wire _09640_;
 wire _09641_;
 wire _09642_;
 wire _09643_;
 wire _09644_;
 wire _09645_;
 wire _09646_;
 wire _09647_;
 wire _09648_;
 wire _09649_;
 wire _09650_;
 wire _09651_;
 wire _09652_;
 wire _09653_;
 wire _09654_;
 wire _09655_;
 wire _09656_;
 wire _09657_;
 wire _09658_;
 wire _09659_;
 wire _09660_;
 wire _09661_;
 wire _09662_;
 wire _09663_;
 wire _09664_;
 wire _09665_;
 wire _09666_;
 wire _09667_;
 wire _09668_;
 wire _09669_;
 wire _09670_;
 wire _09671_;
 wire _09672_;
 wire _09673_;
 wire _09674_;
 wire _09675_;
 wire _09676_;
 wire _09677_;
 wire _09678_;
 wire _09679_;
 wire _09680_;
 wire _09681_;
 wire _09682_;
 wire _09683_;
 wire _09684_;
 wire _09685_;
 wire _09686_;
 wire _09687_;
 wire _09688_;
 wire _09689_;
 wire _09690_;
 wire _09691_;
 wire _09692_;
 wire _09693_;
 wire _09694_;
 wire _09695_;
 wire _09696_;
 wire _09697_;
 wire _09698_;
 wire _09699_;
 wire _09700_;
 wire _09701_;
 wire _09702_;
 wire _09703_;
 wire _09704_;
 wire _09705_;
 wire _09706_;
 wire _09707_;
 wire _09708_;
 wire _09709_;
 wire _09710_;
 wire _09711_;
 wire _09712_;
 wire net610;
 wire _09714_;
 wire net7;
 wire net4;
 wire _09717_;
 wire _09718_;
 wire _09719_;
 wire net138;
 wire net174;
 wire _09722_;
 wire _09723_;
 wire _09724_;
 wire _09725_;
 wire _09726_;
 wire _09727_;
 wire _09728_;
 wire _09729_;
 wire _09730_;
 wire _09731_;
 wire _09732_;
 wire _09733_;
 wire _09734_;
 wire _09735_;
 wire _09736_;
 wire net12;
 wire net145;
 wire _09739_;
 wire _09740_;
 wire _09741_;
 wire _09742_;
 wire _09743_;
 wire _09744_;
 wire _09745_;
 wire _09746_;
 wire _09747_;
 wire _09748_;
 wire _09749_;
 wire _09750_;
 wire _09751_;
 wire _09752_;
 wire _09753_;
 wire _09754_;
 wire _09755_;
 wire _09756_;
 wire net617;
 wire net173;
 wire _09759_;
 wire _09760_;
 wire _09761_;
 wire _09762_;
 wire _09763_;
 wire _09764_;
 wire _09765_;
 wire _09766_;
 wire _09767_;
 wire _09768_;
 wire _09769_;
 wire _09770_;
 wire _09771_;
 wire _09772_;
 wire _09773_;
 wire _09774_;
 wire _09775_;
 wire _09776_;
 wire _09777_;
 wire _09778_;
 wire _09779_;
 wire _09780_;
 wire _09781_;
 wire _09782_;
 wire _09783_;
 wire _09784_;
 wire _09785_;
 wire _09786_;
 wire _09787_;
 wire _09788_;
 wire _09789_;
 wire _09790_;
 wire _09791_;
 wire _09792_;
 wire _09793_;
 wire _09794_;
 wire _09795_;
 wire _09796_;
 wire _09797_;
 wire _09798_;
 wire _09799_;
 wire _09800_;
 wire _09801_;
 wire _09802_;
 wire _09803_;
 wire _09804_;
 wire _09805_;
 wire _09806_;
 wire _09807_;
 wire _09808_;
 wire _09809_;
 wire _09810_;
 wire _09811_;
 wire _09812_;
 wire _09813_;
 wire _09814_;
 wire _09815_;
 wire _09816_;
 wire _09817_;
 wire _09818_;
 wire _09819_;
 wire _09820_;
 wire _09821_;
 wire _09822_;
 wire _09823_;
 wire _09824_;
 wire _09825_;
 wire _09826_;
 wire _09827_;
 wire _09828_;
 wire _09829_;
 wire _09830_;
 wire _09831_;
 wire _09832_;
 wire _09833_;
 wire _09834_;
 wire _09835_;
 wire _09836_;
 wire _09837_;
 wire _09838_;
 wire _09839_;
 wire _09840_;
 wire _09841_;
 wire _09842_;
 wire _09843_;
 wire _09844_;
 wire _09845_;
 wire _09846_;
 wire _09847_;
 wire _09848_;
 wire _09849_;
 wire _09850_;
 wire _09851_;
 wire _09852_;
 wire _09853_;
 wire _09854_;
 wire _09855_;
 wire _09856_;
 wire _09857_;
 wire _09858_;
 wire _09859_;
 wire _09860_;
 wire _09861_;
 wire _09862_;
 wire _09863_;
 wire _09864_;
 wire _09865_;
 wire _09866_;
 wire _09867_;
 wire _09868_;
 wire _09869_;
 wire _09870_;
 wire _09871_;
 wire _09872_;
 wire _09873_;
 wire _09874_;
 wire _09875_;
 wire _09876_;
 wire _09877_;
 wire _09878_;
 wire _09879_;
 wire _09880_;
 wire _09881_;
 wire _09882_;
 wire net160;
 wire _09884_;
 wire _09885_;
 wire _09886_;
 wire _09887_;
 wire _09888_;
 wire _09889_;
 wire _09890_;
 wire _09891_;
 wire _09892_;
 wire _09893_;
 wire _09894_;
 wire _09895_;
 wire _09896_;
 wire _09897_;
 wire _09898_;
 wire net15;
 wire _09900_;
 wire _09901_;
 wire _09902_;
 wire _09903_;
 wire _09904_;
 wire _09905_;
 wire net144;
 wire _09907_;
 wire _09908_;
 wire _09909_;
 wire _09910_;
 wire _09911_;
 wire _09912_;
 wire _09913_;
 wire _09914_;
 wire _09915_;
 wire _09916_;
 wire _09917_;
 wire _09918_;
 wire _09919_;
 wire _09920_;
 wire _09921_;
 wire _09922_;
 wire _09923_;
 wire _09924_;
 wire _09925_;
 wire _09926_;
 wire _09927_;
 wire _09928_;
 wire _09929_;
 wire _09930_;
 wire _09931_;
 wire _09932_;
 wire _09933_;
 wire _09934_;
 wire _09935_;
 wire _09936_;
 wire _09937_;
 wire _09938_;
 wire _09939_;
 wire _09940_;
 wire _09941_;
 wire _09942_;
 wire _09943_;
 wire _09944_;
 wire _09945_;
 wire _09946_;
 wire _09947_;
 wire _09948_;
 wire _09949_;
 wire _09950_;
 wire _09951_;
 wire net107;
 wire _09953_;
 wire _09954_;
 wire _09955_;
 wire _09956_;
 wire _09957_;
 wire _09958_;
 wire _09959_;
 wire _09960_;
 wire _09961_;
 wire _09962_;
 wire _09963_;
 wire _09964_;
 wire _09965_;
 wire _09966_;
 wire _09967_;
 wire _09968_;
 wire _09969_;
 wire _09970_;
 wire _09971_;
 wire _09972_;
 wire _09973_;
 wire _09974_;
 wire _09975_;
 wire _09976_;
 wire _09977_;
 wire _09978_;
 wire _09979_;
 wire _09980_;
 wire _09981_;
 wire _09982_;
 wire _09983_;
 wire _09984_;
 wire _09985_;
 wire _09986_;
 wire _09987_;
 wire _09988_;
 wire _09989_;
 wire _09990_;
 wire _09991_;
 wire _09992_;
 wire _09993_;
 wire _09994_;
 wire _09995_;
 wire _09996_;
 wire _09997_;
 wire _09998_;
 wire _09999_;
 wire _10000_;
 wire _10001_;
 wire _10002_;
 wire _10003_;
 wire _10004_;
 wire _10005_;
 wire _10006_;
 wire _10007_;
 wire _10008_;
 wire _10009_;
 wire _10010_;
 wire _10011_;
 wire _10012_;
 wire _10013_;
 wire _10014_;
 wire _10015_;
 wire _10016_;
 wire _10017_;
 wire _10018_;
 wire _10019_;
 wire _10020_;
 wire _10021_;
 wire _10022_;
 wire _10023_;
 wire _10024_;
 wire _10025_;
 wire _10026_;
 wire _10027_;
 wire _10028_;
 wire _10029_;
 wire _10030_;
 wire _10031_;
 wire _10032_;
 wire _10033_;
 wire _10034_;
 wire _10035_;
 wire _10036_;
 wire _10037_;
 wire _10038_;
 wire _10039_;
 wire _10040_;
 wire _10041_;
 wire _10042_;
 wire _10043_;
 wire _10044_;
 wire _10045_;
 wire _10046_;
 wire _10047_;
 wire _10048_;
 wire _10049_;
 wire _10050_;
 wire _10051_;
 wire _10052_;
 wire _10053_;
 wire _10054_;
 wire _10055_;
 wire _10056_;
 wire _10057_;
 wire _10058_;
 wire _10059_;
 wire _10060_;
 wire _10061_;
 wire _10062_;
 wire _10063_;
 wire _10064_;
 wire _10065_;
 wire _10066_;
 wire _10067_;
 wire _10068_;
 wire _10069_;
 wire _10070_;
 wire _10071_;
 wire _10072_;
 wire _10073_;
 wire _10074_;
 wire _10075_;
 wire _10076_;
 wire _10077_;
 wire _10078_;
 wire _10079_;
 wire _10080_;
 wire _10081_;
 wire _10082_;
 wire _10083_;
 wire _10084_;
 wire _10085_;
 wire _10086_;
 wire _10087_;
 wire _10088_;
 wire _10089_;
 wire _10090_;
 wire _10091_;
 wire _10092_;
 wire _10093_;
 wire _10094_;
 wire _10095_;
 wire _10096_;
 wire _10097_;
 wire _10098_;
 wire _10099_;
 wire _10100_;
 wire _10101_;
 wire _10102_;
 wire _10103_;
 wire _10104_;
 wire _10105_;
 wire _10106_;
 wire _10107_;
 wire _10108_;
 wire _10109_;
 wire _10110_;
 wire _10111_;
 wire _10112_;
 wire _10113_;
 wire _10114_;
 wire _10115_;
 wire _10116_;
 wire _10117_;
 wire _10118_;
 wire _10119_;
 wire _10120_;
 wire _10121_;
 wire _10122_;
 wire _10123_;
 wire _10124_;
 wire _10125_;
 wire _10126_;
 wire _10127_;
 wire _10128_;
 wire _10129_;
 wire _10130_;
 wire _10131_;
 wire _10132_;
 wire _10133_;
 wire _10134_;
 wire _10135_;
 wire _10136_;
 wire _10137_;
 wire _10138_;
 wire _10139_;
 wire _10140_;
 wire _10141_;
 wire _10142_;
 wire _10143_;
 wire _10144_;
 wire _10145_;
 wire _10146_;
 wire _10147_;
 wire _10148_;
 wire _10149_;
 wire _10150_;
 wire _10151_;
 wire _10152_;
 wire _10153_;
 wire _10154_;
 wire _10155_;
 wire _10156_;
 wire _10157_;
 wire _10158_;
 wire _10159_;
 wire _10160_;
 wire _10161_;
 wire _10162_;
 wire _10163_;
 wire _10164_;
 wire _10165_;
 wire _10166_;
 wire _10167_;
 wire _10168_;
 wire _10169_;
 wire _10170_;
 wire _10171_;
 wire _10172_;
 wire _10173_;
 wire _10174_;
 wire _10175_;
 wire _10176_;
 wire _10177_;
 wire _10178_;
 wire _10179_;
 wire _10180_;
 wire _10181_;
 wire _10182_;
 wire _10183_;
 wire _10184_;
 wire _10185_;
 wire _10186_;
 wire _10187_;
 wire _10188_;
 wire _10189_;
 wire _10190_;
 wire _10191_;
 wire _10192_;
 wire _10193_;
 wire _10194_;
 wire _10195_;
 wire _10196_;
 wire _10197_;
 wire _10198_;
 wire _10199_;
 wire _10200_;
 wire _10201_;
 wire _10202_;
 wire _10203_;
 wire _10204_;
 wire _10205_;
 wire _10206_;
 wire _10207_;
 wire _10208_;
 wire _10209_;
 wire _10210_;
 wire _10211_;
 wire _10212_;
 wire _10213_;
 wire _10214_;
 wire _10215_;
 wire _10216_;
 wire _10217_;
 wire _10218_;
 wire _10219_;
 wire _10220_;
 wire _10221_;
 wire _10222_;
 wire _10223_;
 wire _10224_;
 wire _10225_;
 wire _10226_;
 wire _10227_;
 wire _10228_;
 wire _10229_;
 wire _10230_;
 wire _10231_;
 wire _10232_;
 wire _10233_;
 wire _10234_;
 wire _10235_;
 wire _10236_;
 wire _10237_;
 wire _10238_;
 wire _10239_;
 wire _10240_;
 wire _10241_;
 wire _10242_;
 wire _10243_;
 wire _10244_;
 wire _10245_;
 wire _10246_;
 wire _10247_;
 wire _10248_;
 wire _10249_;
 wire _10250_;
 wire _10251_;
 wire _10252_;
 wire _10253_;
 wire _10254_;
 wire _10255_;
 wire _10256_;
 wire _10257_;
 wire _10258_;
 wire _10259_;
 wire _10260_;
 wire _10261_;
 wire _10262_;
 wire _10263_;
 wire _10264_;
 wire _10265_;
 wire _10266_;
 wire _10267_;
 wire _10268_;
 wire _10269_;
 wire _10270_;
 wire _10271_;
 wire _10272_;
 wire _10273_;
 wire _10274_;
 wire _10275_;
 wire _10276_;
 wire _10277_;
 wire _10278_;
 wire _10279_;
 wire _10280_;
 wire _10281_;
 wire _10282_;
 wire _10283_;
 wire _10284_;
 wire _10285_;
 wire _10286_;
 wire _10287_;
 wire _10288_;
 wire _10289_;
 wire _10290_;
 wire _10291_;
 wire _10292_;
 wire _10293_;
 wire _10294_;
 wire _10295_;
 wire _10296_;
 wire _10297_;
 wire _10298_;
 wire _10299_;
 wire _10300_;
 wire _10301_;
 wire _10302_;
 wire _10303_;
 wire _10304_;
 wire _10305_;
 wire _10306_;
 wire _10307_;
 wire _10308_;
 wire _10309_;
 wire _10310_;
 wire _10311_;
 wire _10312_;
 wire _10313_;
 wire _10314_;
 wire _10315_;
 wire _10316_;
 wire _10317_;
 wire _10318_;
 wire _10319_;
 wire _10320_;
 wire _10321_;
 wire _10322_;
 wire _10323_;
 wire _10324_;
 wire _10325_;
 wire _10326_;
 wire _10327_;
 wire _10328_;
 wire _10329_;
 wire _10330_;
 wire _10331_;
 wire _10332_;
 wire _10333_;
 wire _10334_;
 wire _10335_;
 wire _10336_;
 wire _10337_;
 wire _10338_;
 wire _10339_;
 wire _10340_;
 wire _10341_;
 wire _10342_;
 wire _10343_;
 wire _10344_;
 wire _10345_;
 wire _10346_;
 wire _10347_;
 wire _10348_;
 wire _10349_;
 wire _10350_;
 wire _10351_;
 wire _10352_;
 wire _10353_;
 wire _10354_;
 wire _10355_;
 wire _10356_;
 wire _10357_;
 wire _10358_;
 wire _10359_;
 wire _10360_;
 wire _10361_;
 wire _10362_;
 wire _10363_;
 wire _10364_;
 wire _10365_;
 wire _10366_;
 wire _10367_;
 wire _10368_;
 wire _10369_;
 wire _10370_;
 wire _10371_;
 wire _10372_;
 wire _10373_;
 wire _10374_;
 wire _10375_;
 wire _10376_;
 wire _10377_;
 wire _10378_;
 wire _10379_;
 wire _10380_;
 wire _10381_;
 wire _10382_;
 wire _10383_;
 wire _10384_;
 wire _10385_;
 wire _10386_;
 wire _10387_;
 wire _10388_;
 wire _10389_;
 wire _10390_;
 wire _10391_;
 wire _10392_;
 wire _10393_;
 wire _10394_;
 wire _10395_;
 wire _10396_;
 wire _10397_;
 wire _10398_;
 wire _10399_;
 wire _10400_;
 wire _10401_;
 wire _10402_;
 wire _10403_;
 wire _10404_;
 wire _10405_;
 wire _10406_;
 wire _10407_;
 wire _10408_;
 wire _10409_;
 wire _10410_;
 wire _10411_;
 wire _10412_;
 wire _10413_;
 wire _10414_;
 wire _10415_;
 wire _10416_;
 wire _10417_;
 wire _10418_;
 wire _10419_;
 wire _10420_;
 wire _10421_;
 wire _10422_;
 wire _10423_;
 wire _10424_;
 wire _10425_;
 wire _10426_;
 wire _10427_;
 wire _10428_;
 wire _10429_;
 wire _10430_;
 wire _10431_;
 wire _10432_;
 wire net537;
 wire _10434_;
 wire net95;
 wire net96;
 wire _10437_;
 wire _10438_;
 wire _10439_;
 wire net5;
 wire net153;
 wire _10442_;
 wire _10443_;
 wire _10444_;
 wire _10445_;
 wire _10446_;
 wire _10447_;
 wire _10448_;
 wire _10449_;
 wire _10450_;
 wire _10451_;
 wire _10452_;
 wire _10453_;
 wire net57;
 wire _10455_;
 wire _10456_;
 wire _10457_;
 wire _10458_;
 wire _10459_;
 wire _10460_;
 wire _10461_;
 wire _10462_;
 wire _10463_;
 wire _10464_;
 wire _10465_;
 wire _10466_;
 wire _10467_;
 wire _10468_;
 wire _10469_;
 wire _10470_;
 wire _10471_;
 wire _10472_;
 wire _10473_;
 wire net133;
 wire _10475_;
 wire _10476_;
 wire _10477_;
 wire _10478_;
 wire _10479_;
 wire _10480_;
 wire _10481_;
 wire _10482_;
 wire _10483_;
 wire _10484_;
 wire _10485_;
 wire _10486_;
 wire _10487_;
 wire _10488_;
 wire _10489_;
 wire _10490_;
 wire _10491_;
 wire _10492_;
 wire _10493_;
 wire _10494_;
 wire _10495_;
 wire _10496_;
 wire _10497_;
 wire _10498_;
 wire _10499_;
 wire _10500_;
 wire _10501_;
 wire _10502_;
 wire _10503_;
 wire _10504_;
 wire _10505_;
 wire _10506_;
 wire _10507_;
 wire _10508_;
 wire _10509_;
 wire _10510_;
 wire _10511_;
 wire _10512_;
 wire _10513_;
 wire _10514_;
 wire _10515_;
 wire _10516_;
 wire _10517_;
 wire _10518_;
 wire _10519_;
 wire _10520_;
 wire _10521_;
 wire _10522_;
 wire _10523_;
 wire _10524_;
 wire _10525_;
 wire _10526_;
 wire _10527_;
 wire _10528_;
 wire _10529_;
 wire _10530_;
 wire _10531_;
 wire _10532_;
 wire _10533_;
 wire _10534_;
 wire _10535_;
 wire _10536_;
 wire _10537_;
 wire _10538_;
 wire _10539_;
 wire _10540_;
 wire _10541_;
 wire _10542_;
 wire _10543_;
 wire _10544_;
 wire _10545_;
 wire _10546_;
 wire _10547_;
 wire _10548_;
 wire _10549_;
 wire _10550_;
 wire _10551_;
 wire _10552_;
 wire _10553_;
 wire _10554_;
 wire _10555_;
 wire _10556_;
 wire _10557_;
 wire _10558_;
 wire _10559_;
 wire _10560_;
 wire _10561_;
 wire _10562_;
 wire _10563_;
 wire _10564_;
 wire _10565_;
 wire _10566_;
 wire _10567_;
 wire _10568_;
 wire _10569_;
 wire _10570_;
 wire _10571_;
 wire _10572_;
 wire _10573_;
 wire _10574_;
 wire _10575_;
 wire _10576_;
 wire _10577_;
 wire _10578_;
 wire _10579_;
 wire _10580_;
 wire _10581_;
 wire _10582_;
 wire _10583_;
 wire _10584_;
 wire _10585_;
 wire _10586_;
 wire _10587_;
 wire _10588_;
 wire _10589_;
 wire _10590_;
 wire _10591_;
 wire _10592_;
 wire _10593_;
 wire _10594_;
 wire _10595_;
 wire _10596_;
 wire _10597_;
 wire _10598_;
 wire _10599_;
 wire _10600_;
 wire _10601_;
 wire _10602_;
 wire _10603_;
 wire _10604_;
 wire _10605_;
 wire _10606_;
 wire _10607_;
 wire net165;
 wire _10609_;
 wire _10610_;
 wire _10611_;
 wire _10612_;
 wire _10613_;
 wire _10614_;
 wire _10615_;
 wire _10616_;
 wire _10617_;
 wire _10618_;
 wire _10619_;
 wire _10620_;
 wire _10621_;
 wire _10622_;
 wire _10623_;
 wire _10624_;
 wire _10625_;
 wire _10626_;
 wire _10627_;
 wire _10628_;
 wire _10629_;
 wire _10630_;
 wire _10631_;
 wire _10632_;
 wire _10633_;
 wire _10634_;
 wire _10635_;
 wire _10636_;
 wire _10637_;
 wire _10638_;
 wire _10639_;
 wire _10640_;
 wire _10641_;
 wire _10642_;
 wire _10643_;
 wire _10644_;
 wire _10645_;
 wire _10646_;
 wire _10647_;
 wire _10648_;
 wire _10649_;
 wire _10650_;
 wire _10651_;
 wire _10652_;
 wire _10653_;
 wire _10654_;
 wire _10655_;
 wire _10656_;
 wire _10657_;
 wire _10658_;
 wire _10659_;
 wire _10660_;
 wire _10661_;
 wire _10662_;
 wire _10663_;
 wire _10664_;
 wire _10665_;
 wire _10666_;
 wire _10667_;
 wire _10668_;
 wire _10669_;
 wire _10670_;
 wire _10671_;
 wire _10672_;
 wire _10673_;
 wire _10674_;
 wire _10675_;
 wire net152;
 wire _10677_;
 wire _10678_;
 wire _10679_;
 wire _10680_;
 wire _10681_;
 wire _10682_;
 wire _10683_;
 wire _10684_;
 wire _10685_;
 wire _10686_;
 wire _10687_;
 wire _10688_;
 wire _10689_;
 wire _10690_;
 wire _10691_;
 wire _10692_;
 wire _10693_;
 wire _10694_;
 wire _10695_;
 wire _10696_;
 wire _10697_;
 wire _10698_;
 wire _10699_;
 wire _10700_;
 wire _10701_;
 wire _10702_;
 wire _10703_;
 wire _10704_;
 wire _10705_;
 wire _10706_;
 wire _10707_;
 wire _10708_;
 wire _10709_;
 wire _10710_;
 wire _10711_;
 wire _10712_;
 wire _10713_;
 wire _10714_;
 wire _10715_;
 wire _10716_;
 wire _10717_;
 wire _10718_;
 wire _10719_;
 wire _10720_;
 wire _10721_;
 wire _10722_;
 wire _10723_;
 wire _10724_;
 wire _10725_;
 wire _10726_;
 wire _10727_;
 wire _10728_;
 wire _10729_;
 wire _10730_;
 wire _10731_;
 wire _10732_;
 wire _10733_;
 wire _10734_;
 wire _10735_;
 wire _10736_;
 wire _10737_;
 wire _10738_;
 wire _10739_;
 wire _10740_;
 wire _10741_;
 wire _10742_;
 wire _10743_;
 wire _10744_;
 wire _10745_;
 wire _10746_;
 wire _10747_;
 wire _10748_;
 wire _10749_;
 wire _10750_;
 wire _10751_;
 wire _10752_;
 wire _10753_;
 wire _10754_;
 wire _10755_;
 wire _10756_;
 wire _10757_;
 wire _10758_;
 wire _10759_;
 wire _10760_;
 wire _10761_;
 wire _10762_;
 wire _10763_;
 wire _10764_;
 wire _10765_;
 wire _10766_;
 wire _10767_;
 wire _10768_;
 wire _10769_;
 wire _10770_;
 wire _10771_;
 wire _10772_;
 wire _10773_;
 wire _10774_;
 wire _10775_;
 wire _10776_;
 wire _10777_;
 wire _10778_;
 wire _10779_;
 wire _10780_;
 wire _10781_;
 wire _10782_;
 wire _10783_;
 wire _10784_;
 wire _10785_;
 wire _10786_;
 wire _10787_;
 wire _10788_;
 wire _10789_;
 wire _10790_;
 wire _10791_;
 wire _10792_;
 wire _10793_;
 wire _10794_;
 wire _10795_;
 wire _10796_;
 wire _10797_;
 wire _10798_;
 wire _10799_;
 wire _10800_;
 wire _10801_;
 wire _10802_;
 wire _10803_;
 wire _10804_;
 wire _10805_;
 wire _10806_;
 wire _10807_;
 wire _10808_;
 wire _10809_;
 wire _10810_;
 wire _10811_;
 wire _10812_;
 wire _10813_;
 wire _10814_;
 wire _10815_;
 wire _10816_;
 wire _10817_;
 wire _10818_;
 wire _10819_;
 wire _10820_;
 wire _10821_;
 wire _10822_;
 wire _10823_;
 wire _10824_;
 wire _10825_;
 wire _10826_;
 wire _10827_;
 wire _10828_;
 wire _10829_;
 wire _10830_;
 wire _10831_;
 wire _10832_;
 wire _10833_;
 wire _10834_;
 wire _10835_;
 wire _10836_;
 wire _10837_;
 wire _10838_;
 wire _10839_;
 wire _10840_;
 wire _10841_;
 wire _10842_;
 wire _10843_;
 wire _10844_;
 wire _10845_;
 wire _10846_;
 wire _10847_;
 wire _10848_;
 wire _10849_;
 wire _10850_;
 wire _10851_;
 wire _10852_;
 wire _10853_;
 wire _10854_;
 wire _10855_;
 wire _10856_;
 wire _10857_;
 wire _10858_;
 wire _10859_;
 wire _10860_;
 wire _10861_;
 wire _10862_;
 wire _10863_;
 wire _10864_;
 wire _10865_;
 wire _10866_;
 wire _10867_;
 wire _10868_;
 wire _10869_;
 wire _10870_;
 wire _10871_;
 wire _10872_;
 wire _10873_;
 wire _10874_;
 wire _10875_;
 wire _10876_;
 wire _10877_;
 wire _10878_;
 wire _10879_;
 wire _10880_;
 wire _10881_;
 wire _10882_;
 wire _10883_;
 wire _10884_;
 wire _10885_;
 wire _10886_;
 wire _10887_;
 wire _10888_;
 wire _10889_;
 wire _10890_;
 wire _10891_;
 wire _10892_;
 wire _10893_;
 wire _10894_;
 wire _10895_;
 wire _10896_;
 wire _10897_;
 wire _10898_;
 wire _10899_;
 wire _10900_;
 wire _10901_;
 wire _10902_;
 wire _10903_;
 wire _10904_;
 wire _10905_;
 wire _10906_;
 wire _10907_;
 wire _10908_;
 wire _10909_;
 wire _10910_;
 wire _10911_;
 wire _10912_;
 wire _10913_;
 wire _10914_;
 wire _10915_;
 wire _10916_;
 wire _10917_;
 wire _10918_;
 wire _10919_;
 wire _10920_;
 wire _10921_;
 wire _10922_;
 wire _10923_;
 wire _10924_;
 wire _10925_;
 wire _10926_;
 wire _10927_;
 wire _10928_;
 wire _10929_;
 wire _10930_;
 wire _10931_;
 wire _10932_;
 wire _10933_;
 wire _10934_;
 wire _10935_;
 wire _10936_;
 wire _10937_;
 wire _10938_;
 wire _10939_;
 wire _10940_;
 wire _10941_;
 wire _10942_;
 wire _10943_;
 wire _10944_;
 wire _10945_;
 wire _10946_;
 wire _10947_;
 wire _10948_;
 wire _10949_;
 wire _10950_;
 wire _10951_;
 wire _10952_;
 wire _10953_;
 wire _10954_;
 wire _10955_;
 wire _10956_;
 wire _10957_;
 wire _10958_;
 wire _10959_;
 wire _10960_;
 wire _10961_;
 wire _10962_;
 wire _10963_;
 wire _10964_;
 wire _10965_;
 wire _10966_;
 wire _10967_;
 wire _10968_;
 wire _10969_;
 wire _10970_;
 wire _10971_;
 wire _10972_;
 wire _10973_;
 wire _10974_;
 wire _10975_;
 wire _10976_;
 wire _10977_;
 wire _10978_;
 wire _10979_;
 wire _10980_;
 wire _10981_;
 wire _10982_;
 wire _10983_;
 wire _10984_;
 wire _10985_;
 wire _10986_;
 wire _10987_;
 wire _10988_;
 wire _10989_;
 wire _10990_;
 wire _10991_;
 wire _10992_;
 wire _10993_;
 wire _10994_;
 wire _10995_;
 wire _10996_;
 wire _10997_;
 wire _10998_;
 wire _10999_;
 wire _11000_;
 wire _11001_;
 wire _11002_;
 wire _11003_;
 wire _11004_;
 wire _11005_;
 wire _11006_;
 wire _11007_;
 wire _11008_;
 wire _11009_;
 wire _11010_;
 wire _11011_;
 wire _11012_;
 wire _11013_;
 wire _11014_;
 wire _11015_;
 wire _11016_;
 wire _11017_;
 wire _11018_;
 wire _11019_;
 wire _11020_;
 wire _11021_;
 wire _11022_;
 wire _11023_;
 wire _11024_;
 wire _11025_;
 wire _11026_;
 wire _11027_;
 wire _11028_;
 wire _11029_;
 wire _11030_;
 wire _11031_;
 wire _11032_;
 wire _11033_;
 wire _11034_;
 wire _11035_;
 wire _11036_;
 wire _11037_;
 wire _11038_;
 wire _11039_;
 wire _11040_;
 wire _11041_;
 wire _11042_;
 wire _11043_;
 wire _11044_;
 wire _11045_;
 wire _11046_;
 wire _11047_;
 wire _11048_;
 wire _11049_;
 wire _11050_;
 wire _11051_;
 wire _11052_;
 wire _11053_;
 wire _11054_;
 wire _11055_;
 wire _11056_;
 wire _11057_;
 wire _11058_;
 wire _11059_;
 wire _11060_;
 wire _11061_;
 wire _11062_;
 wire _11063_;
 wire _11064_;
 wire _11065_;
 wire _11066_;
 wire _11067_;
 wire _11068_;
 wire _11069_;
 wire _11070_;
 wire _11071_;
 wire _11072_;
 wire _11073_;
 wire _11074_;
 wire _11075_;
 wire _11076_;
 wire _11077_;
 wire _11078_;
 wire _11079_;
 wire _11080_;
 wire _11081_;
 wire _11082_;
 wire _11083_;
 wire _11084_;
 wire _11085_;
 wire _11086_;
 wire _11087_;
 wire _11088_;
 wire _11089_;
 wire _11090_;
 wire _11091_;
 wire _11092_;
 wire _11093_;
 wire _11094_;
 wire _11095_;
 wire _11096_;
 wire _11097_;
 wire _11098_;
 wire _11099_;
 wire _11100_;
 wire _11101_;
 wire _11102_;
 wire _11103_;
 wire _11104_;
 wire _11105_;
 wire _11106_;
 wire _11107_;
 wire _11108_;
 wire _11109_;
 wire _11110_;
 wire _11111_;
 wire _11112_;
 wire _11113_;
 wire _11114_;
 wire net102;
 wire net65;
 wire _11117_;
 wire _11118_;
 wire _11119_;
 wire _11120_;
 wire _11121_;
 wire _11122_;
 wire _11123_;
 wire _11124_;
 wire _11125_;
 wire _11126_;
 wire _11127_;
 wire _11128_;
 wire _11129_;
 wire _11130_;
 wire _11131_;
 wire net590;
 wire _11133_;
 wire _11134_;
 wire _11135_;
 wire _11136_;
 wire _11137_;
 wire _11138_;
 wire _11139_;
 wire _11140_;
 wire _11141_;
 wire _11142_;
 wire _11143_;
 wire _11144_;
 wire _11145_;
 wire _11146_;
 wire _11147_;
 wire _11148_;
 wire _11149_;
 wire _11150_;
 wire _11151_;
 wire _11152_;
 wire _11153_;
 wire _11154_;
 wire _11155_;
 wire _11156_;
 wire _11157_;
 wire _11158_;
 wire _11159_;
 wire _11160_;
 wire _11161_;
 wire _11162_;
 wire _11163_;
 wire _11164_;
 wire net657;
 wire _11166_;
 wire _11167_;
 wire _11168_;
 wire _11169_;
 wire _11170_;
 wire _11171_;
 wire _11172_;
 wire _11173_;
 wire _11174_;
 wire _11175_;
 wire _11176_;
 wire _11177_;
 wire _11178_;
 wire _11179_;
 wire _11180_;
 wire _11181_;
 wire _11182_;
 wire _11183_;
 wire _11184_;
 wire _11185_;
 wire _11186_;
 wire _11187_;
 wire _11188_;
 wire _11189_;
 wire _11190_;
 wire _11191_;
 wire _11192_;
 wire _11193_;
 wire _11194_;
 wire _11195_;
 wire _11196_;
 wire _11197_;
 wire _11198_;
 wire _11199_;
 wire _11200_;
 wire _11201_;
 wire _11202_;
 wire _11203_;
 wire _11204_;
 wire _11205_;
 wire _11206_;
 wire _11207_;
 wire _11208_;
 wire _11209_;
 wire _11210_;
 wire _11211_;
 wire _11212_;
 wire net49;
 wire _11214_;
 wire _11215_;
 wire _11216_;
 wire _11217_;
 wire _11218_;
 wire _11219_;
 wire _11220_;
 wire _11221_;
 wire _11222_;
 wire _11223_;
 wire _11224_;
 wire _11225_;
 wire _11226_;
 wire _11227_;
 wire _11228_;
 wire _11229_;
 wire _11230_;
 wire _11231_;
 wire _11232_;
 wire _11233_;
 wire _11234_;
 wire _11235_;
 wire _11236_;
 wire _11237_;
 wire _11238_;
 wire _11239_;
 wire _11240_;
 wire _11241_;
 wire _11242_;
 wire _11243_;
 wire _11244_;
 wire _11245_;
 wire _11246_;
 wire _11247_;
 wire _11248_;
 wire _11249_;
 wire _11250_;
 wire _11251_;
 wire _11252_;
 wire _11253_;
 wire _11254_;
 wire _11255_;
 wire _11256_;
 wire _11257_;
 wire _11258_;
 wire _11259_;
 wire _11260_;
 wire _11261_;
 wire _11262_;
 wire _11263_;
 wire _11264_;
 wire _11265_;
 wire _11266_;
 wire _11267_;
 wire _11268_;
 wire _11269_;
 wire _11270_;
 wire _11271_;
 wire _11272_;
 wire _11273_;
 wire _11274_;
 wire _11275_;
 wire _11276_;
 wire _11277_;
 wire _11278_;
 wire _11279_;
 wire _11280_;
 wire _11281_;
 wire _11282_;
 wire _11283_;
 wire _11284_;
 wire _11285_;
 wire _11286_;
 wire _11287_;
 wire _11288_;
 wire _11289_;
 wire _11290_;
 wire _11291_;
 wire _11292_;
 wire _11293_;
 wire _11294_;
 wire _11295_;
 wire _11296_;
 wire _11297_;
 wire _11298_;
 wire _11299_;
 wire _11300_;
 wire _11301_;
 wire net9;
 wire _11303_;
 wire _11304_;
 wire _11305_;
 wire _11306_;
 wire _11307_;
 wire _11308_;
 wire _11309_;
 wire _11310_;
 wire net43;
 wire _11312_;
 wire _11313_;
 wire _11314_;
 wire _11315_;
 wire _11316_;
 wire _11317_;
 wire _11318_;
 wire _11319_;
 wire _11320_;
 wire _11321_;
 wire _11322_;
 wire _11323_;
 wire _11324_;
 wire _11325_;
 wire _11326_;
 wire _11327_;
 wire _11328_;
 wire _11329_;
 wire _11330_;
 wire _11331_;
 wire _11332_;
 wire _11333_;
 wire _11334_;
 wire _11335_;
 wire _11336_;
 wire _11337_;
 wire _11338_;
 wire _11339_;
 wire _11340_;
 wire _11341_;
 wire _11342_;
 wire _11343_;
 wire _11344_;
 wire _11345_;
 wire _11346_;
 wire _11347_;
 wire _11348_;
 wire _11349_;
 wire _11350_;
 wire _11351_;
 wire _11352_;
 wire _11353_;
 wire _11354_;
 wire _11355_;
 wire _11356_;
 wire _11357_;
 wire _11358_;
 wire _11359_;
 wire _11360_;
 wire _11361_;
 wire _11362_;
 wire _11363_;
 wire _11364_;
 wire _11365_;
 wire _11366_;
 wire _11367_;
 wire _11368_;
 wire _11369_;
 wire _11370_;
 wire _11371_;
 wire _11372_;
 wire _11373_;
 wire _11374_;
 wire _11375_;
 wire _11376_;
 wire _11377_;
 wire _11378_;
 wire _11379_;
 wire _11380_;
 wire _11381_;
 wire _11382_;
 wire _11383_;
 wire _11384_;
 wire _11385_;
 wire _11386_;
 wire _11387_;
 wire _11388_;
 wire _11389_;
 wire _11390_;
 wire _11391_;
 wire _11392_;
 wire _11393_;
 wire _11394_;
 wire _11395_;
 wire _11396_;
 wire _11397_;
 wire _11398_;
 wire _11399_;
 wire _11400_;
 wire _11401_;
 wire _11402_;
 wire _11403_;
 wire _11404_;
 wire _11405_;
 wire _11406_;
 wire _11407_;
 wire _11408_;
 wire _11409_;
 wire _11410_;
 wire _11411_;
 wire _11412_;
 wire _11413_;
 wire _11414_;
 wire _11415_;
 wire _11416_;
 wire _11417_;
 wire _11418_;
 wire _11419_;
 wire _11420_;
 wire _11421_;
 wire _11422_;
 wire _11423_;
 wire _11424_;
 wire _11425_;
 wire _11426_;
 wire _11427_;
 wire _11428_;
 wire _11429_;
 wire _11430_;
 wire _11431_;
 wire _11432_;
 wire _11433_;
 wire _11434_;
 wire _11435_;
 wire _11436_;
 wire _11437_;
 wire _11438_;
 wire _11439_;
 wire _11440_;
 wire _11441_;
 wire _11442_;
 wire _11443_;
 wire _11444_;
 wire _11445_;
 wire _11446_;
 wire _11447_;
 wire _11448_;
 wire _11449_;
 wire _11450_;
 wire _11451_;
 wire _11452_;
 wire _11453_;
 wire _11454_;
 wire _11455_;
 wire _11456_;
 wire _11457_;
 wire _11458_;
 wire _11459_;
 wire _11460_;
 wire _11461_;
 wire _11462_;
 wire _11463_;
 wire _11464_;
 wire _11465_;
 wire _11466_;
 wire _11467_;
 wire _11468_;
 wire _11469_;
 wire _11470_;
 wire _11471_;
 wire _11472_;
 wire _11473_;
 wire _11474_;
 wire _11475_;
 wire _11476_;
 wire _11477_;
 wire _11478_;
 wire _11479_;
 wire _11480_;
 wire _11481_;
 wire _11482_;
 wire _11483_;
 wire _11484_;
 wire _11485_;
 wire _11486_;
 wire _11487_;
 wire _11488_;
 wire _11489_;
 wire _11490_;
 wire _11491_;
 wire _11492_;
 wire _11493_;
 wire _11494_;
 wire _11495_;
 wire _11496_;
 wire _11497_;
 wire _11498_;
 wire _11499_;
 wire _11500_;
 wire _11501_;
 wire _11502_;
 wire _11503_;
 wire _11504_;
 wire _11505_;
 wire _11506_;
 wire _11507_;
 wire _11508_;
 wire _11509_;
 wire _11510_;
 wire _11511_;
 wire _11512_;
 wire _11513_;
 wire _11514_;
 wire _11515_;
 wire _11516_;
 wire _11517_;
 wire _11518_;
 wire _11519_;
 wire _11520_;
 wire _11521_;
 wire _11522_;
 wire _11523_;
 wire _11524_;
 wire _11525_;
 wire _11526_;
 wire _11527_;
 wire _11528_;
 wire _11529_;
 wire _11530_;
 wire _11531_;
 wire _11532_;
 wire _11533_;
 wire _11534_;
 wire _11535_;
 wire _11536_;
 wire _11537_;
 wire _11538_;
 wire _11539_;
 wire _11540_;
 wire _11541_;
 wire _11542_;
 wire _11543_;
 wire _11544_;
 wire _11545_;
 wire _11546_;
 wire _11547_;
 wire _11548_;
 wire _11549_;
 wire _11550_;
 wire _11551_;
 wire _11552_;
 wire _11553_;
 wire _11554_;
 wire _11555_;
 wire _11556_;
 wire _11557_;
 wire _11558_;
 wire _11559_;
 wire _11560_;
 wire _11561_;
 wire _11562_;
 wire _11563_;
 wire _11564_;
 wire _11565_;
 wire _11566_;
 wire _11567_;
 wire _11568_;
 wire _11569_;
 wire _11570_;
 wire _11571_;
 wire _11572_;
 wire _11573_;
 wire _11574_;
 wire _11575_;
 wire _11576_;
 wire _11577_;
 wire _11578_;
 wire _11579_;
 wire _11580_;
 wire _11581_;
 wire _11582_;
 wire _11583_;
 wire _11584_;
 wire _11585_;
 wire _11586_;
 wire _11587_;
 wire _11588_;
 wire _11589_;
 wire _11590_;
 wire _11591_;
 wire _11592_;
 wire _11593_;
 wire _11594_;
 wire _11595_;
 wire _11596_;
 wire _11597_;
 wire _11598_;
 wire _11599_;
 wire _11600_;
 wire _11601_;
 wire _11602_;
 wire _11603_;
 wire _11604_;
 wire _11605_;
 wire _11606_;
 wire _11607_;
 wire _11608_;
 wire _11609_;
 wire _11610_;
 wire _11611_;
 wire _11612_;
 wire _11613_;
 wire _11614_;
 wire _11615_;
 wire _11616_;
 wire _11617_;
 wire _11618_;
 wire _11619_;
 wire _11620_;
 wire _11621_;
 wire _11622_;
 wire _11623_;
 wire _11624_;
 wire _11625_;
 wire _11626_;
 wire _11627_;
 wire _11628_;
 wire _11629_;
 wire _11630_;
 wire _11631_;
 wire _11632_;
 wire _11633_;
 wire _11634_;
 wire _11635_;
 wire _11636_;
 wire _11637_;
 wire _11638_;
 wire _11639_;
 wire _11640_;
 wire _11641_;
 wire _11642_;
 wire _11643_;
 wire _11644_;
 wire _11645_;
 wire _11646_;
 wire _11647_;
 wire _11648_;
 wire _11649_;
 wire _11650_;
 wire _11651_;
 wire _11652_;
 wire _11653_;
 wire _11654_;
 wire _11655_;
 wire _11656_;
 wire _11657_;
 wire _11658_;
 wire _11659_;
 wire _11660_;
 wire _11661_;
 wire _11662_;
 wire _11663_;
 wire _11664_;
 wire _11665_;
 wire _11666_;
 wire _11667_;
 wire _11668_;
 wire _11669_;
 wire _11670_;
 wire _11671_;
 wire _11672_;
 wire _11673_;
 wire _11674_;
 wire _11675_;
 wire _11676_;
 wire _11677_;
 wire _11678_;
 wire _11679_;
 wire _11680_;
 wire _11681_;
 wire _11682_;
 wire _11683_;
 wire _11684_;
 wire _11685_;
 wire _11686_;
 wire _11687_;
 wire _11688_;
 wire _11689_;
 wire _11690_;
 wire _11691_;
 wire _11692_;
 wire _11693_;
 wire _11694_;
 wire _11695_;
 wire _11696_;
 wire _11697_;
 wire _11698_;
 wire _11699_;
 wire _11700_;
 wire _11701_;
 wire _11702_;
 wire _11703_;
 wire _11704_;
 wire _11705_;
 wire _11706_;
 wire _11707_;
 wire _11708_;
 wire _11709_;
 wire _11710_;
 wire _11711_;
 wire _11712_;
 wire _11713_;
 wire _11714_;
 wire _11715_;
 wire _11716_;
 wire _11717_;
 wire _11718_;
 wire _11719_;
 wire _11720_;
 wire _11721_;
 wire _11722_;
 wire _11723_;
 wire _11724_;
 wire _11725_;
 wire _11726_;
 wire _11727_;
 wire _11728_;
 wire _11729_;
 wire _11730_;
 wire _11731_;
 wire _11732_;
 wire _11733_;
 wire _11734_;
 wire _11735_;
 wire _11736_;
 wire _11737_;
 wire _11738_;
 wire _11739_;
 wire _11740_;
 wire _11741_;
 wire _11742_;
 wire _11743_;
 wire _11744_;
 wire _11745_;
 wire _11746_;
 wire _11747_;
 wire _11748_;
 wire _11749_;
 wire _11750_;
 wire _11751_;
 wire _11752_;
 wire _11753_;
 wire _11754_;
 wire _11755_;
 wire _11756_;
 wire _11757_;
 wire _11758_;
 wire _11759_;
 wire _11760_;
 wire _11761_;
 wire _11762_;
 wire _11763_;
 wire _11764_;
 wire _11765_;
 wire _11766_;
 wire _11767_;
 wire _11768_;
 wire _11769_;
 wire _11770_;
 wire _11771_;
 wire _11772_;
 wire _11773_;
 wire _11774_;
 wire _11775_;
 wire _11776_;
 wire _11777_;
 wire _11778_;
 wire _11779_;
 wire _11780_;
 wire _11781_;
 wire _11782_;
 wire _11783_;
 wire _11784_;
 wire _11785_;
 wire _11786_;
 wire _11787_;
 wire _11788_;
 wire _11789_;
 wire _11790_;
 wire _11791_;
 wire _11792_;
 wire _11793_;
 wire _11794_;
 wire _11795_;
 wire _11796_;
 wire _11797_;
 wire _11798_;
 wire _11799_;
 wire _11800_;
 wire _11801_;
 wire _11802_;
 wire _11803_;
 wire _11804_;
 wire _11805_;
 wire _11806_;
 wire _11807_;
 wire _11808_;
 wire _11809_;
 wire _11810_;
 wire _11811_;
 wire _11812_;
 wire _11813_;
 wire _11814_;
 wire _11815_;
 wire _11816_;
 wire _11817_;
 wire _11818_;
 wire _11819_;
 wire _11820_;
 wire _11821_;
 wire _11822_;
 wire _11823_;
 wire _11824_;
 wire _11825_;
 wire _11826_;
 wire _11827_;
 wire _11828_;
 wire _11829_;
 wire _11830_;
 wire _11831_;
 wire _11832_;
 wire _11833_;
 wire _11834_;
 wire _11835_;
 wire _11836_;
 wire _11837_;
 wire _11838_;
 wire _11839_;
 wire _11840_;
 wire _11841_;
 wire _11842_;
 wire _11843_;
 wire _11844_;
 wire _11845_;
 wire _11846_;
 wire _11847_;
 wire _11848_;
 wire _11849_;
 wire _11850_;
 wire _11851_;
 wire _11852_;
 wire _11853_;
 wire net109;
 wire _11855_;
 wire _11856_;
 wire _11857_;
 wire _11858_;
 wire _11859_;
 wire _11860_;
 wire _11861_;
 wire _11862_;
 wire _11863_;
 wire _11864_;
 wire _11865_;
 wire _11866_;
 wire _11867_;
 wire _11868_;
 wire _11869_;
 wire _11870_;
 wire _11871_;
 wire _11872_;
 wire _11873_;
 wire _11874_;
 wire _11875_;
 wire _11876_;
 wire _11877_;
 wire _11878_;
 wire _11879_;
 wire _11880_;
 wire _11881_;
 wire _11882_;
 wire _11883_;
 wire _11884_;
 wire _11885_;
 wire _11886_;
 wire _11887_;
 wire _11888_;
 wire _11889_;
 wire _11890_;
 wire _11891_;
 wire _11892_;
 wire _11893_;
 wire _11894_;
 wire _11895_;
 wire _11896_;
 wire _11897_;
 wire _11898_;
 wire _11899_;
 wire _11900_;
 wire _11901_;
 wire _11902_;
 wire _11903_;
 wire _11904_;
 wire _11905_;
 wire _11906_;
 wire _11907_;
 wire _11908_;
 wire _11909_;
 wire _11910_;
 wire _11911_;
 wire _11912_;
 wire _11913_;
 wire _11914_;
 wire _11915_;
 wire _11916_;
 wire _11917_;
 wire _11918_;
 wire _11919_;
 wire _11920_;
 wire _11921_;
 wire _11922_;
 wire _11923_;
 wire _11924_;
 wire _11925_;
 wire _11926_;
 wire _11927_;
 wire _11928_;
 wire _11929_;
 wire _11930_;
 wire _11931_;
 wire _11932_;
 wire _11933_;
 wire _11934_;
 wire net110;
 wire _11936_;
 wire _11937_;
 wire _11938_;
 wire _11939_;
 wire _11940_;
 wire _11941_;
 wire _11942_;
 wire _11943_;
 wire _11944_;
 wire _11945_;
 wire _11946_;
 wire _11947_;
 wire _11948_;
 wire _11949_;
 wire _11950_;
 wire _11951_;
 wire _11952_;
 wire _11953_;
 wire _11954_;
 wire _11955_;
 wire _11956_;
 wire _11957_;
 wire _11958_;
 wire _11959_;
 wire _11960_;
 wire _11961_;
 wire _11962_;
 wire _11963_;
 wire _11964_;
 wire _11965_;
 wire _11966_;
 wire _11967_;
 wire _11968_;
 wire _11969_;
 wire _11970_;
 wire _11971_;
 wire _11972_;
 wire _11973_;
 wire _11974_;
 wire _11975_;
 wire _11976_;
 wire _11977_;
 wire _11978_;
 wire _11979_;
 wire _11980_;
 wire _11981_;
 wire _11982_;
 wire _11983_;
 wire _11984_;
 wire _11985_;
 wire _11986_;
 wire _11987_;
 wire _11988_;
 wire _11989_;
 wire _11990_;
 wire _11991_;
 wire _11992_;
 wire _11993_;
 wire _11994_;
 wire _11995_;
 wire _11996_;
 wire _11997_;
 wire _11998_;
 wire _11999_;
 wire _12000_;
 wire _12001_;
 wire _12002_;
 wire _12003_;
 wire _12004_;
 wire _12005_;
 wire _12006_;
 wire _12007_;
 wire _12008_;
 wire _12009_;
 wire _12010_;
 wire _12011_;
 wire _12012_;
 wire _12013_;
 wire _12014_;
 wire _12015_;
 wire _12016_;
 wire _12017_;
 wire _12018_;
 wire _12019_;
 wire _12020_;
 wire _12021_;
 wire _12022_;
 wire _12023_;
 wire _12024_;
 wire _12025_;
 wire _12026_;
 wire _12027_;
 wire _12028_;
 wire _12029_;
 wire _12030_;
 wire _12031_;
 wire _12032_;
 wire _12033_;
 wire _12034_;
 wire _12035_;
 wire _12036_;
 wire _12037_;
 wire _12038_;
 wire _12039_;
 wire _12040_;
 wire _12041_;
 wire _12042_;
 wire _12043_;
 wire _12044_;
 wire _12045_;
 wire _12046_;
 wire _12047_;
 wire net1098;
 wire _12049_;
 wire _12050_;
 wire _12051_;
 wire _12052_;
 wire _12053_;
 wire _12054_;
 wire _12055_;
 wire _12056_;
 wire _12057_;
 wire _12058_;
 wire _12059_;
 wire _12060_;
 wire _12061_;
 wire _12062_;
 wire _12063_;
 wire _12064_;
 wire _12065_;
 wire _12066_;
 wire _12067_;
 wire _12068_;
 wire _12069_;
 wire _12070_;
 wire _12071_;
 wire _12072_;
 wire _12073_;
 wire _12074_;
 wire _12075_;
 wire _12076_;
 wire _12077_;
 wire _12078_;
 wire _12079_;
 wire _12080_;
 wire _12081_;
 wire _12082_;
 wire _12083_;
 wire _12084_;
 wire _12085_;
 wire _12086_;
 wire _12087_;
 wire _12088_;
 wire _12089_;
 wire _12090_;
 wire _12091_;
 wire _12092_;
 wire _12093_;
 wire _12094_;
 wire _12095_;
 wire _12096_;
 wire _12097_;
 wire _12098_;
 wire _12099_;
 wire _12100_;
 wire _12101_;
 wire _12102_;
 wire _12103_;
 wire _12104_;
 wire _12105_;
 wire _12106_;
 wire _12107_;
 wire _12108_;
 wire _12109_;
 wire _12110_;
 wire _12111_;
 wire _12112_;
 wire _12113_;
 wire _12114_;
 wire _12115_;
 wire _12116_;
 wire _12117_;
 wire _12118_;
 wire _12119_;
 wire _12120_;
 wire _12121_;
 wire _12122_;
 wire _12123_;
 wire _12124_;
 wire _12125_;
 wire _12126_;
 wire _12127_;
 wire _12128_;
 wire _12129_;
 wire _12130_;
 wire _12131_;
 wire _12132_;
 wire _12133_;
 wire _12134_;
 wire _12135_;
 wire _12136_;
 wire _12137_;
 wire _12138_;
 wire _12139_;
 wire _12140_;
 wire _12141_;
 wire _12142_;
 wire _12143_;
 wire _12144_;
 wire _12145_;
 wire _12146_;
 wire _12147_;
 wire _12148_;
 wire _12149_;
 wire _12150_;
 wire _12151_;
 wire _12152_;
 wire _12153_;
 wire _12154_;
 wire _12155_;
 wire _12156_;
 wire _12157_;
 wire _12158_;
 wire _12159_;
 wire _12160_;
 wire _12161_;
 wire _12162_;
 wire _12163_;
 wire _12164_;
 wire _12165_;
 wire _12166_;
 wire _12167_;
 wire _12168_;
 wire _12169_;
 wire _12170_;
 wire _12171_;
 wire _12172_;
 wire _12173_;
 wire _12174_;
 wire _12175_;
 wire _12176_;
 wire _12177_;
 wire _12178_;
 wire _12179_;
 wire _12180_;
 wire _12181_;
 wire _12182_;
 wire _12183_;
 wire _12184_;
 wire _12185_;
 wire _12186_;
 wire _12187_;
 wire _12188_;
 wire _12189_;
 wire _12190_;
 wire _12191_;
 wire _12192_;
 wire _12193_;
 wire _12194_;
 wire _12195_;
 wire _12196_;
 wire _12197_;
 wire _12198_;
 wire _12199_;
 wire _12200_;
 wire _12201_;
 wire _12202_;
 wire _12203_;
 wire _12204_;
 wire _12205_;
 wire _12206_;
 wire _12207_;
 wire _12208_;
 wire _12209_;
 wire _12210_;
 wire _12211_;
 wire _12212_;
 wire _12213_;
 wire _12214_;
 wire _12215_;
 wire _12216_;
 wire _12217_;
 wire _12218_;
 wire _12219_;
 wire _12220_;
 wire _12221_;
 wire _12222_;
 wire _12223_;
 wire _12224_;
 wire _12225_;
 wire _12226_;
 wire _12227_;
 wire _12228_;
 wire _12229_;
 wire _12230_;
 wire _12231_;
 wire _12232_;
 wire _12233_;
 wire _12234_;
 wire _12235_;
 wire _12236_;
 wire _12237_;
 wire _12238_;
 wire _12239_;
 wire _12240_;
 wire _12241_;
 wire _12242_;
 wire _12243_;
 wire _12244_;
 wire _12245_;
 wire _12246_;
 wire _12247_;
 wire _12248_;
 wire _12249_;
 wire _12250_;
 wire _12251_;
 wire _12252_;
 wire _12253_;
 wire _12254_;
 wire _12255_;
 wire _12256_;
 wire _12257_;
 wire _12258_;
 wire _12259_;
 wire _12260_;
 wire _12261_;
 wire _12262_;
 wire _12263_;
 wire _12264_;
 wire _12265_;
 wire _12266_;
 wire _12267_;
 wire _12268_;
 wire _12269_;
 wire _12270_;
 wire _12271_;
 wire _12272_;
 wire _12273_;
 wire _12274_;
 wire _12275_;
 wire _12276_;
 wire _12277_;
 wire _12278_;
 wire _12279_;
 wire _12280_;
 wire _12281_;
 wire _12282_;
 wire _12283_;
 wire _12284_;
 wire _12285_;
 wire _12286_;
 wire _12287_;
 wire _12288_;
 wire _12289_;
 wire _12290_;
 wire _12291_;
 wire _12292_;
 wire _12293_;
 wire _12294_;
 wire _12295_;
 wire _12296_;
 wire _12297_;
 wire _12298_;
 wire _12299_;
 wire _12300_;
 wire _12301_;
 wire _12302_;
 wire _12303_;
 wire _12304_;
 wire _12305_;
 wire _12306_;
 wire _12307_;
 wire _12308_;
 wire _12309_;
 wire _12310_;
 wire _12311_;
 wire _12312_;
 wire _12313_;
 wire _12314_;
 wire _12315_;
 wire _12316_;
 wire _12317_;
 wire _12318_;
 wire _12319_;
 wire _12320_;
 wire _12321_;
 wire _12322_;
 wire _12323_;
 wire _12324_;
 wire _12325_;
 wire _12326_;
 wire _12327_;
 wire _12328_;
 wire _12329_;
 wire _12330_;
 wire _12331_;
 wire _12332_;
 wire _12333_;
 wire _12334_;
 wire _12335_;
 wire _12336_;
 wire _12337_;
 wire _12338_;
 wire _12339_;
 wire _12340_;
 wire _12341_;
 wire _12342_;
 wire _12343_;
 wire _12344_;
 wire _12345_;
 wire _12346_;
 wire _12347_;
 wire _12348_;
 wire _12349_;
 wire _12350_;
 wire _12351_;
 wire _12352_;
 wire _12353_;
 wire _12354_;
 wire _12355_;
 wire _12356_;
 wire _12357_;
 wire _12358_;
 wire _12359_;
 wire _12360_;
 wire _12361_;
 wire _12362_;
 wire _12363_;
 wire _12364_;
 wire _12365_;
 wire _12366_;
 wire _12367_;
 wire _12368_;
 wire _12369_;
 wire _12370_;
 wire _12371_;
 wire _12372_;
 wire _12373_;
 wire _12374_;
 wire _12375_;
 wire _12376_;
 wire _12377_;
 wire _12378_;
 wire _12379_;
 wire _12380_;
 wire _12381_;
 wire _12382_;
 wire _12383_;
 wire _12384_;
 wire _12385_;
 wire _12386_;
 wire _12387_;
 wire _12388_;
 wire _12389_;
 wire _12390_;
 wire _12391_;
 wire _12392_;
 wire _12393_;
 wire _12394_;
 wire _12395_;
 wire _12396_;
 wire _12397_;
 wire _12398_;
 wire _12399_;
 wire _12400_;
 wire _12401_;
 wire _12402_;
 wire _12403_;
 wire _12404_;
 wire _12405_;
 wire _12406_;
 wire _12407_;
 wire _12408_;
 wire _12409_;
 wire _12410_;
 wire _12411_;
 wire _12412_;
 wire _12413_;
 wire _12414_;
 wire _12415_;
 wire _12416_;
 wire _12417_;
 wire _12418_;
 wire _12419_;
 wire _12420_;
 wire _12421_;
 wire _12422_;
 wire _12423_;
 wire _12424_;
 wire _12425_;
 wire _12426_;
 wire _12427_;
 wire _12428_;
 wire _12429_;
 wire _12430_;
 wire _12431_;
 wire _12432_;
 wire _12433_;
 wire _12434_;
 wire _12435_;
 wire _12436_;
 wire _12437_;
 wire _12438_;
 wire _12439_;
 wire _12440_;
 wire _12441_;
 wire _12442_;
 wire _12443_;
 wire _12444_;
 wire _12445_;
 wire _12446_;
 wire _12447_;
 wire _12448_;
 wire _12449_;
 wire _12450_;
 wire _12451_;
 wire _12452_;
 wire _12453_;
 wire _12454_;
 wire _12455_;
 wire _12456_;
 wire _12457_;
 wire _12458_;
 wire _12459_;
 wire _12460_;
 wire _12461_;
 wire _12462_;
 wire _12463_;
 wire _12464_;
 wire _12465_;
 wire _12466_;
 wire _12467_;
 wire _12468_;
 wire _12469_;
 wire _12470_;
 wire _12471_;
 wire _12472_;
 wire _12473_;
 wire _12474_;
 wire _12475_;
 wire _12476_;
 wire _12477_;
 wire _12478_;
 wire _12479_;
 wire _12480_;
 wire _12481_;
 wire _12482_;
 wire _12483_;
 wire _12484_;
 wire _12485_;
 wire _12486_;
 wire _12487_;
 wire _12488_;
 wire _12489_;
 wire _12490_;
 wire _12491_;
 wire _12492_;
 wire _12493_;
 wire _12494_;
 wire _12495_;
 wire _12496_;
 wire _12497_;
 wire _12498_;
 wire _12499_;
 wire _12500_;
 wire _12501_;
 wire _12502_;
 wire _12503_;
 wire _12504_;
 wire _12505_;
 wire _12506_;
 wire net139;
 wire _12508_;
 wire net1162;
 wire _12510_;
 wire _12511_;
 wire _12512_;
 wire _12513_;
 wire _12514_;
 wire _12515_;
 wire _12516_;
 wire _12517_;
 wire _12518_;
 wire _12519_;
 wire _12520_;
 wire _12521_;
 wire _12522_;
 wire _12523_;
 wire _12524_;
 wire _12525_;
 wire _12526_;
 wire _12527_;
 wire net98;
 wire _12529_;
 wire _12530_;
 wire _12531_;
 wire _12532_;
 wire _12533_;
 wire _12534_;
 wire _12535_;
 wire _12536_;
 wire _12537_;
 wire _12538_;
 wire _12539_;
 wire _12540_;
 wire _12541_;
 wire _12542_;
 wire _12543_;
 wire _12544_;
 wire _12545_;
 wire _12546_;
 wire _12547_;
 wire _12548_;
 wire _12549_;
 wire _12550_;
 wire _12551_;
 wire _12552_;
 wire _12553_;
 wire _12554_;
 wire _12555_;
 wire _12556_;
 wire _12557_;
 wire _12558_;
 wire _12559_;
 wire _12560_;
 wire _12561_;
 wire _12562_;
 wire _12563_;
 wire _12564_;
 wire _12565_;
 wire _12566_;
 wire _12567_;
 wire _12568_;
 wire _12569_;
 wire _12570_;
 wire _12571_;
 wire _12572_;
 wire _12573_;
 wire _12574_;
 wire _12575_;
 wire _12576_;
 wire _12577_;
 wire _12578_;
 wire _12579_;
 wire _12580_;
 wire _12581_;
 wire _12582_;
 wire _12583_;
 wire _12584_;
 wire net146;
 wire _12586_;
 wire _12587_;
 wire _12588_;
 wire _12589_;
 wire _12590_;
 wire _12591_;
 wire _12592_;
 wire _12593_;
 wire _12594_;
 wire _12595_;
 wire _12596_;
 wire _12597_;
 wire _12598_;
 wire _12599_;
 wire _12600_;
 wire _12601_;
 wire _12602_;
 wire _12603_;
 wire _12604_;
 wire _12605_;
 wire _12606_;
 wire _12607_;
 wire _12608_;
 wire _12609_;
 wire _12610_;
 wire _12611_;
 wire _12612_;
 wire _12613_;
 wire _12614_;
 wire _12615_;
 wire _12616_;
 wire _12617_;
 wire _12618_;
 wire _12619_;
 wire _12620_;
 wire _12621_;
 wire _12622_;
 wire _12623_;
 wire _12624_;
 wire _12625_;
 wire _12626_;
 wire _12627_;
 wire _12628_;
 wire _12629_;
 wire _12630_;
 wire _12631_;
 wire _12632_;
 wire _12633_;
 wire _12634_;
 wire _12635_;
 wire _12636_;
 wire _12637_;
 wire _12638_;
 wire _12639_;
 wire _12640_;
 wire net166;
 wire _12642_;
 wire _12643_;
 wire _12644_;
 wire _12645_;
 wire _12646_;
 wire _12647_;
 wire net140;
 wire _12649_;
 wire _12650_;
 wire _12651_;
 wire _12652_;
 wire net171;
 wire _12654_;
 wire _12655_;
 wire _12656_;
 wire _12657_;
 wire _12658_;
 wire _12659_;
 wire _12660_;
 wire _12661_;
 wire _12662_;
 wire _12663_;
 wire _12664_;
 wire _12665_;
 wire _12666_;
 wire _12667_;
 wire _12668_;
 wire _12669_;
 wire _12670_;
 wire net914;
 wire _12672_;
 wire _12673_;
 wire _12674_;
 wire _12675_;
 wire _12676_;
 wire _12677_;
 wire _12678_;
 wire _12679_;
 wire _12680_;
 wire _12681_;
 wire _12682_;
 wire _12683_;
 wire _12684_;
 wire _12685_;
 wire _12686_;
 wire _12687_;
 wire _12688_;
 wire _12689_;
 wire _12690_;
 wire _12691_;
 wire _12692_;
 wire _12693_;
 wire _12694_;
 wire _12695_;
 wire _12696_;
 wire _12697_;
 wire _12698_;
 wire _12699_;
 wire _12700_;
 wire _12701_;
 wire _12702_;
 wire _12703_;
 wire _12704_;
 wire _12705_;
 wire _12706_;
 wire _12707_;
 wire _12708_;
 wire _12709_;
 wire _12710_;
 wire _12711_;
 wire _12712_;
 wire _12713_;
 wire _12714_;
 wire _12715_;
 wire _12716_;
 wire _12717_;
 wire _12718_;
 wire _12719_;
 wire _12720_;
 wire _12721_;
 wire _12722_;
 wire _12723_;
 wire _12724_;
 wire _12725_;
 wire _12726_;
 wire _12727_;
 wire _12728_;
 wire _12729_;
 wire _12730_;
 wire _12731_;
 wire _12732_;
 wire _12733_;
 wire _12734_;
 wire _12735_;
 wire _12736_;
 wire _12737_;
 wire _12738_;
 wire _12739_;
 wire _12740_;
 wire _12741_;
 wire _12742_;
 wire _12743_;
 wire _12744_;
 wire _12745_;
 wire _12746_;
 wire _12747_;
 wire _12748_;
 wire _12749_;
 wire _12750_;
 wire _12751_;
 wire _12752_;
 wire _12753_;
 wire _12754_;
 wire _12755_;
 wire _12756_;
 wire _12757_;
 wire _12758_;
 wire _12759_;
 wire _12760_;
 wire _12761_;
 wire _12762_;
 wire _12763_;
 wire _12764_;
 wire _12765_;
 wire _12766_;
 wire _12767_;
 wire _12768_;
 wire _12769_;
 wire _12770_;
 wire _12771_;
 wire _12772_;
 wire _12773_;
 wire _12774_;
 wire _12775_;
 wire _12776_;
 wire _12777_;
 wire _12778_;
 wire _12779_;
 wire _12780_;
 wire _12781_;
 wire _12782_;
 wire _12783_;
 wire _12784_;
 wire _12785_;
 wire _12786_;
 wire _12787_;
 wire _12788_;
 wire _12789_;
 wire _12790_;
 wire _12791_;
 wire _12792_;
 wire _12793_;
 wire _12794_;
 wire _12795_;
 wire _12796_;
 wire _12797_;
 wire _12798_;
 wire _12799_;
 wire _12800_;
 wire _12801_;
 wire _12802_;
 wire _12803_;
 wire _12804_;
 wire _12805_;
 wire _12806_;
 wire _12807_;
 wire _12808_;
 wire _12809_;
 wire _12810_;
 wire _12811_;
 wire _12812_;
 wire _12813_;
 wire _12814_;
 wire _12815_;
 wire _12816_;
 wire _12817_;
 wire _12818_;
 wire _12819_;
 wire _12820_;
 wire _12821_;
 wire _12822_;
 wire _12823_;
 wire _12824_;
 wire _12825_;
 wire _12826_;
 wire _12827_;
 wire _12828_;
 wire _12829_;
 wire _12830_;
 wire _12831_;
 wire _12832_;
 wire _12833_;
 wire _12834_;
 wire _12835_;
 wire _12836_;
 wire _12837_;
 wire _12838_;
 wire _12839_;
 wire _12840_;
 wire _12841_;
 wire _12842_;
 wire _12843_;
 wire _12844_;
 wire _12845_;
 wire _12846_;
 wire _12847_;
 wire _12848_;
 wire _12849_;
 wire _12850_;
 wire _12851_;
 wire _12852_;
 wire _12853_;
 wire _12854_;
 wire _12855_;
 wire _12856_;
 wire _12857_;
 wire _12858_;
 wire _12859_;
 wire _12860_;
 wire _12861_;
 wire _12862_;
 wire _12863_;
 wire _12864_;
 wire _12865_;
 wire _12866_;
 wire _12867_;
 wire _12868_;
 wire _12869_;
 wire _12870_;
 wire _12871_;
 wire _12872_;
 wire _12873_;
 wire _12874_;
 wire _12875_;
 wire _12876_;
 wire _12877_;
 wire _12878_;
 wire _12879_;
 wire _12880_;
 wire _12881_;
 wire _12882_;
 wire _12883_;
 wire _12884_;
 wire _12885_;
 wire _12886_;
 wire _12887_;
 wire _12888_;
 wire _12889_;
 wire _12890_;
 wire _12891_;
 wire _12892_;
 wire _12893_;
 wire _12894_;
 wire _12895_;
 wire _12896_;
 wire _12897_;
 wire _12898_;
 wire _12899_;
 wire _12900_;
 wire _12901_;
 wire _12902_;
 wire _12903_;
 wire _12904_;
 wire _12905_;
 wire _12906_;
 wire _12907_;
 wire _12908_;
 wire _12909_;
 wire _12910_;
 wire _12911_;
 wire _12912_;
 wire _12913_;
 wire _12914_;
 wire _12915_;
 wire _12916_;
 wire _12917_;
 wire _12918_;
 wire _12919_;
 wire _12920_;
 wire _12921_;
 wire _12922_;
 wire _12923_;
 wire _12924_;
 wire _12925_;
 wire _12926_;
 wire _12927_;
 wire _12928_;
 wire _12929_;
 wire _12930_;
 wire _12931_;
 wire _12932_;
 wire _12933_;
 wire _12934_;
 wire _12935_;
 wire _12936_;
 wire _12937_;
 wire _12938_;
 wire _12939_;
 wire _12940_;
 wire _12941_;
 wire _12942_;
 wire _12943_;
 wire _12944_;
 wire _12945_;
 wire _12946_;
 wire _12947_;
 wire _12948_;
 wire _12949_;
 wire _12950_;
 wire _12951_;
 wire _12952_;
 wire _12953_;
 wire _12954_;
 wire _12955_;
 wire _12956_;
 wire _12957_;
 wire _12958_;
 wire _12959_;
 wire _12960_;
 wire _12961_;
 wire _12962_;
 wire _12963_;
 wire _12964_;
 wire _12965_;
 wire _12966_;
 wire _12967_;
 wire _12968_;
 wire _12969_;
 wire _12970_;
 wire _12971_;
 wire _12972_;
 wire _12973_;
 wire _12974_;
 wire _12975_;
 wire _12976_;
 wire _12977_;
 wire _12978_;
 wire _12979_;
 wire _12980_;
 wire _12981_;
 wire _12982_;
 wire _12983_;
 wire _12984_;
 wire _12985_;
 wire _12986_;
 wire _12987_;
 wire _12988_;
 wire _12989_;
 wire _12990_;
 wire _12991_;
 wire _12992_;
 wire _12993_;
 wire _12994_;
 wire _12995_;
 wire _12996_;
 wire _12997_;
 wire _12998_;
 wire _12999_;
 wire _13000_;
 wire _13001_;
 wire _13002_;
 wire _13003_;
 wire _13004_;
 wire _13005_;
 wire _13006_;
 wire _13007_;
 wire _13008_;
 wire _13009_;
 wire _13010_;
 wire _13011_;
 wire _13012_;
 wire _13013_;
 wire _13014_;
 wire _13015_;
 wire _13016_;
 wire _13017_;
 wire _13018_;
 wire _13019_;
 wire _13020_;
 wire _13021_;
 wire _13022_;
 wire _13023_;
 wire _13024_;
 wire _13025_;
 wire _13026_;
 wire _13027_;
 wire _13028_;
 wire _13029_;
 wire _13030_;
 wire _13031_;
 wire _13032_;
 wire _13033_;
 wire _13034_;
 wire _13035_;
 wire _13036_;
 wire _13037_;
 wire _13038_;
 wire _13039_;
 wire _13040_;
 wire _13041_;
 wire _13042_;
 wire _13043_;
 wire _13044_;
 wire _13045_;
 wire _13046_;
 wire _13047_;
 wire _13048_;
 wire _13049_;
 wire _13050_;
 wire _13051_;
 wire _13052_;
 wire _13053_;
 wire _13054_;
 wire _13055_;
 wire _13056_;
 wire _13057_;
 wire _13058_;
 wire _13059_;
 wire _13060_;
 wire _13061_;
 wire _13062_;
 wire _13063_;
 wire _13064_;
 wire _13065_;
 wire _13066_;
 wire _13067_;
 wire _13068_;
 wire _13069_;
 wire _13070_;
 wire _13071_;
 wire _13072_;
 wire _13073_;
 wire _13074_;
 wire _13075_;
 wire _13076_;
 wire _13077_;
 wire _13078_;
 wire _13079_;
 wire _13080_;
 wire _13081_;
 wire _13082_;
 wire _13083_;
 wire _13084_;
 wire _13085_;
 wire _13086_;
 wire _13087_;
 wire _13088_;
 wire _13089_;
 wire _13090_;
 wire _13091_;
 wire _13092_;
 wire _13093_;
 wire _13094_;
 wire _13095_;
 wire _13096_;
 wire _13097_;
 wire _13098_;
 wire _13099_;
 wire _13100_;
 wire _13101_;
 wire _13102_;
 wire _13103_;
 wire _13104_;
 wire _13105_;
 wire _13106_;
 wire _13107_;
 wire _13108_;
 wire _13109_;
 wire _13110_;
 wire _13111_;
 wire _13112_;
 wire _13113_;
 wire _13114_;
 wire _13115_;
 wire _13116_;
 wire _13117_;
 wire _13118_;
 wire _13119_;
 wire _13120_;
 wire _13121_;
 wire _13122_;
 wire _13123_;
 wire _13124_;
 wire _13125_;
 wire _13126_;
 wire _13127_;
 wire _13128_;
 wire _13129_;
 wire _13130_;
 wire _13131_;
 wire _13132_;
 wire _13133_;
 wire _13134_;
 wire _13135_;
 wire _13136_;
 wire _13137_;
 wire _13138_;
 wire _13139_;
 wire _13140_;
 wire _13141_;
 wire _13142_;
 wire _13143_;
 wire _13144_;
 wire _13145_;
 wire _13146_;
 wire _13147_;
 wire _13148_;
 wire _13149_;
 wire _13150_;
 wire _13151_;
 wire _13152_;
 wire _13153_;
 wire _13154_;
 wire _13155_;
 wire _13156_;
 wire _13157_;
 wire _13158_;
 wire _13159_;
 wire _13160_;
 wire _13161_;
 wire _13162_;
 wire _13163_;
 wire _13164_;
 wire _13165_;
 wire _13166_;
 wire _13167_;
 wire _13168_;
 wire _13169_;
 wire _13170_;
 wire _13171_;
 wire _13172_;
 wire _13173_;
 wire _13174_;
 wire _13175_;
 wire _13176_;
 wire _13177_;
 wire _13178_;
 wire _13179_;
 wire _13180_;
 wire _13181_;
 wire _13182_;
 wire _13183_;
 wire _13184_;
 wire _13185_;
 wire _13186_;
 wire _13187_;
 wire _13188_;
 wire _13189_;
 wire _13190_;
 wire _13191_;
 wire _13192_;
 wire _13193_;
 wire _13194_;
 wire _13195_;
 wire _13196_;
 wire _13197_;
 wire _13198_;
 wire _13199_;
 wire _13200_;
 wire _13201_;
 wire _13202_;
 wire _13203_;
 wire _13204_;
 wire _13205_;
 wire _13206_;
 wire _13207_;
 wire _13208_;
 wire _13209_;
 wire _13210_;
 wire _13211_;
 wire _13212_;
 wire _13213_;
 wire _13214_;
 wire _13215_;
 wire _13216_;
 wire _13217_;
 wire _13218_;
 wire _13219_;
 wire _13220_;
 wire _13221_;
 wire _13222_;
 wire _13223_;
 wire _13224_;
 wire _13225_;
 wire _13226_;
 wire _13227_;
 wire _13228_;
 wire _13229_;
 wire _13230_;
 wire _13231_;
 wire _13232_;
 wire _13233_;
 wire _13234_;
 wire _13235_;
 wire _13236_;
 wire _13237_;
 wire _13238_;
 wire net141;
 wire _13240_;
 wire _13241_;
 wire _13242_;
 wire _13243_;
 wire _13244_;
 wire _13245_;
 wire _13246_;
 wire _13247_;
 wire _13248_;
 wire _13249_;
 wire _13250_;
 wire _13251_;
 wire _13252_;
 wire _13253_;
 wire _13254_;
 wire _13255_;
 wire _13256_;
 wire _13257_;
 wire _13258_;
 wire _13259_;
 wire _13260_;
 wire _13261_;
 wire _13262_;
 wire _13263_;
 wire _13264_;
 wire _13265_;
 wire _13266_;
 wire _13267_;
 wire _13268_;
 wire _13269_;
 wire _13270_;
 wire _13271_;
 wire _13272_;
 wire _13273_;
 wire _13274_;
 wire _13275_;
 wire _13276_;
 wire _13277_;
 wire _13278_;
 wire _13279_;
 wire _13280_;
 wire _13281_;
 wire _13282_;
 wire _13283_;
 wire _13284_;
 wire _13285_;
 wire _13286_;
 wire _13287_;
 wire _13288_;
 wire _13289_;
 wire _13290_;
 wire _13291_;
 wire _13292_;
 wire _13293_;
 wire _13294_;
 wire _13295_;
 wire _13296_;
 wire _13297_;
 wire _13298_;
 wire _13299_;
 wire _13300_;
 wire _13301_;
 wire _13302_;
 wire _13303_;
 wire _13304_;
 wire _13305_;
 wire _13306_;
 wire _13307_;
 wire _13308_;
 wire _13309_;
 wire _13310_;
 wire _13311_;
 wire net143;
 wire _13313_;
 wire _13314_;
 wire _13315_;
 wire _13316_;
 wire _13317_;
 wire net189;
 wire _13319_;
 wire _13320_;
 wire _13321_;
 wire _13322_;
 wire _13323_;
 wire _13324_;
 wire _13325_;
 wire _13326_;
 wire _13327_;
 wire _13328_;
 wire _13329_;
 wire _13330_;
 wire _13331_;
 wire _13332_;
 wire _13333_;
 wire _13334_;
 wire _13335_;
 wire _13336_;
 wire _13337_;
 wire _13338_;
 wire _13339_;
 wire _13340_;
 wire _13341_;
 wire _13342_;
 wire _13343_;
 wire _13344_;
 wire _13345_;
 wire _13346_;
 wire _13347_;
 wire _13348_;
 wire _13349_;
 wire _13350_;
 wire _13351_;
 wire _13352_;
 wire _13353_;
 wire _13354_;
 wire _13355_;
 wire _13356_;
 wire _13357_;
 wire _13358_;
 wire _13359_;
 wire _13360_;
 wire _13361_;
 wire _13362_;
 wire _13363_;
 wire _13364_;
 wire _13365_;
 wire _13366_;
 wire _13367_;
 wire _13368_;
 wire _13369_;
 wire _13370_;
 wire _13371_;
 wire _13372_;
 wire _13373_;
 wire _13374_;
 wire _13375_;
 wire _13376_;
 wire _13377_;
 wire _13378_;
 wire _13379_;
 wire _13380_;
 wire _13381_;
 wire _13382_;
 wire _13383_;
 wire _13384_;
 wire _13385_;
 wire _13386_;
 wire _13387_;
 wire net632;
 wire _13389_;
 wire _13390_;
 wire _13391_;
 wire _13392_;
 wire _13393_;
 wire _13394_;
 wire _13395_;
 wire _13396_;
 wire _13397_;
 wire _13398_;
 wire _13399_;
 wire _13400_;
 wire _13401_;
 wire _13402_;
 wire _13403_;
 wire _13404_;
 wire _13405_;
 wire _13406_;
 wire _13407_;
 wire _13408_;
 wire _13409_;
 wire _13410_;
 wire _13411_;
 wire _13412_;
 wire _13413_;
 wire _13414_;
 wire _13415_;
 wire _13416_;
 wire _13417_;
 wire _13418_;
 wire _13419_;
 wire _13420_;
 wire _13421_;
 wire _13422_;
 wire _13423_;
 wire _13424_;
 wire _13425_;
 wire _13426_;
 wire _13427_;
 wire _13428_;
 wire _13429_;
 wire _13430_;
 wire _13431_;
 wire _13432_;
 wire _13433_;
 wire _13434_;
 wire _13435_;
 wire _13436_;
 wire _13437_;
 wire _13438_;
 wire _13439_;
 wire _13440_;
 wire _13441_;
 wire _13442_;
 wire _13443_;
 wire _13444_;
 wire _13445_;
 wire _13446_;
 wire _13447_;
 wire _13448_;
 wire _13449_;
 wire _13450_;
 wire _13451_;
 wire _13452_;
 wire _13453_;
 wire _13454_;
 wire _13455_;
 wire _13456_;
 wire _13457_;
 wire _13458_;
 wire _13459_;
 wire _13460_;
 wire _13461_;
 wire _13462_;
 wire _13463_;
 wire _13464_;
 wire _13465_;
 wire _13466_;
 wire _13467_;
 wire _13468_;
 wire _13469_;
 wire _13470_;
 wire _13471_;
 wire _13472_;
 wire _13473_;
 wire _13474_;
 wire _13475_;
 wire _13476_;
 wire _13477_;
 wire _13478_;
 wire _13479_;
 wire _13480_;
 wire _13481_;
 wire _13482_;
 wire _13483_;
 wire _13484_;
 wire _13485_;
 wire _13486_;
 wire _13487_;
 wire _13488_;
 wire _13489_;
 wire _13490_;
 wire _13491_;
 wire _13492_;
 wire _13493_;
 wire _13494_;
 wire _13495_;
 wire _13496_;
 wire _13497_;
 wire _13498_;
 wire _13499_;
 wire _13500_;
 wire _13501_;
 wire _13502_;
 wire _13503_;
 wire _13504_;
 wire _13505_;
 wire _13506_;
 wire _13507_;
 wire _13508_;
 wire _13509_;
 wire _13510_;
 wire _13511_;
 wire _13512_;
 wire _13513_;
 wire _13514_;
 wire _13515_;
 wire _13516_;
 wire _13517_;
 wire _13518_;
 wire _13519_;
 wire _13520_;
 wire _13521_;
 wire _13522_;
 wire _13523_;
 wire _13524_;
 wire _13525_;
 wire _13526_;
 wire _13527_;
 wire _13528_;
 wire _13529_;
 wire _13530_;
 wire _13531_;
 wire _13532_;
 wire _13533_;
 wire _13534_;
 wire _13535_;
 wire _13536_;
 wire _13537_;
 wire _13538_;
 wire _13539_;
 wire _13540_;
 wire _13541_;
 wire _13542_;
 wire _13543_;
 wire _13544_;
 wire _13545_;
 wire _13546_;
 wire _13547_;
 wire _13548_;
 wire _13549_;
 wire _13550_;
 wire _13551_;
 wire _13552_;
 wire _13553_;
 wire _13554_;
 wire _13555_;
 wire _13556_;
 wire _13557_;
 wire _13558_;
 wire _13559_;
 wire _13560_;
 wire _13561_;
 wire _13562_;
 wire _13563_;
 wire _13564_;
 wire _13565_;
 wire _13566_;
 wire _13567_;
 wire _13568_;
 wire _13569_;
 wire _13570_;
 wire _13571_;
 wire _13572_;
 wire _13573_;
 wire _13574_;
 wire _13575_;
 wire _13576_;
 wire _13577_;
 wire _13578_;
 wire _13579_;
 wire _13580_;
 wire _13581_;
 wire _13582_;
 wire _13583_;
 wire _13584_;
 wire _13585_;
 wire _13586_;
 wire _13587_;
 wire _13588_;
 wire _13589_;
 wire _13590_;
 wire _13591_;
 wire _13592_;
 wire _13593_;
 wire _13594_;
 wire _13595_;
 wire _13596_;
 wire _13597_;
 wire _13598_;
 wire _13599_;
 wire _13600_;
 wire _13601_;
 wire _13602_;
 wire _13603_;
 wire _13604_;
 wire _13605_;
 wire _13606_;
 wire _13607_;
 wire _13608_;
 wire _13609_;
 wire _13610_;
 wire _13611_;
 wire _13612_;
 wire _13613_;
 wire _13614_;
 wire _13615_;
 wire _13616_;
 wire _13617_;
 wire _13618_;
 wire _13619_;
 wire _13620_;
 wire _13621_;
 wire _13622_;
 wire _13623_;
 wire _13624_;
 wire _13625_;
 wire _13626_;
 wire _13627_;
 wire _13628_;
 wire _13629_;
 wire _13630_;
 wire _13631_;
 wire _13632_;
 wire _13633_;
 wire _13634_;
 wire _13635_;
 wire _13636_;
 wire _13637_;
 wire _13638_;
 wire _13639_;
 wire _13640_;
 wire _13641_;
 wire _13642_;
 wire _13643_;
 wire _13644_;
 wire _13645_;
 wire _13646_;
 wire _13647_;
 wire _13648_;
 wire _13649_;
 wire _13650_;
 wire _13651_;
 wire _13652_;
 wire _13653_;
 wire _13654_;
 wire _13655_;
 wire _13656_;
 wire _13657_;
 wire _13658_;
 wire _13659_;
 wire _13660_;
 wire _13661_;
 wire _13662_;
 wire _13663_;
 wire _13664_;
 wire _13665_;
 wire _13666_;
 wire _13667_;
 wire _13668_;
 wire _13669_;
 wire _13670_;
 wire _13671_;
 wire _13672_;
 wire _13673_;
 wire _13674_;
 wire _13675_;
 wire _13676_;
 wire _13677_;
 wire _13678_;
 wire _13679_;
 wire _13680_;
 wire _13681_;
 wire _13682_;
 wire _13683_;
 wire _13684_;
 wire _13685_;
 wire _13686_;
 wire _13687_;
 wire _13688_;
 wire _13689_;
 wire _13690_;
 wire _13691_;
 wire _13692_;
 wire _13693_;
 wire _13694_;
 wire _13695_;
 wire _13696_;
 wire _13697_;
 wire _13698_;
 wire _13699_;
 wire _13700_;
 wire _13701_;
 wire _13702_;
 wire _13703_;
 wire _13704_;
 wire _13705_;
 wire _13706_;
 wire _13707_;
 wire _13708_;
 wire _13709_;
 wire _13710_;
 wire _13711_;
 wire _13712_;
 wire _13713_;
 wire _13714_;
 wire _13715_;
 wire _13716_;
 wire _13717_;
 wire _13718_;
 wire _13719_;
 wire _13720_;
 wire _13721_;
 wire _13722_;
 wire _13723_;
 wire _13724_;
 wire _13725_;
 wire _13726_;
 wire _13727_;
 wire _13728_;
 wire _13729_;
 wire _13730_;
 wire _13731_;
 wire _13732_;
 wire _13733_;
 wire _13734_;
 wire _13735_;
 wire _13736_;
 wire _13737_;
 wire _13738_;
 wire _13739_;
 wire _13740_;
 wire _13741_;
 wire _13742_;
 wire _13743_;
 wire _13744_;
 wire _13745_;
 wire _13746_;
 wire _13747_;
 wire _13748_;
 wire _13749_;
 wire _13750_;
 wire _13751_;
 wire _13752_;
 wire _13753_;
 wire _13754_;
 wire _13755_;
 wire _13756_;
 wire _13757_;
 wire _13758_;
 wire _13759_;
 wire _13760_;
 wire _13761_;
 wire _13762_;
 wire _13763_;
 wire _13764_;
 wire _13765_;
 wire _13766_;
 wire _13767_;
 wire _13768_;
 wire _13769_;
 wire _13770_;
 wire _13771_;
 wire _13772_;
 wire _13773_;
 wire _13774_;
 wire _13775_;
 wire _13776_;
 wire _13777_;
 wire _13778_;
 wire _13779_;
 wire _13780_;
 wire _13781_;
 wire _13782_;
 wire _13783_;
 wire _13784_;
 wire _13785_;
 wire _13786_;
 wire _13787_;
 wire _13788_;
 wire _13789_;
 wire _13790_;
 wire _13791_;
 wire _13792_;
 wire _13793_;
 wire _13794_;
 wire _13795_;
 wire _13796_;
 wire _13797_;
 wire _13798_;
 wire _13799_;
 wire _13800_;
 wire _13801_;
 wire _13802_;
 wire _13803_;
 wire _13804_;
 wire _13805_;
 wire _13806_;
 wire _13807_;
 wire _13808_;
 wire _13809_;
 wire _13810_;
 wire _13811_;
 wire _13812_;
 wire _13813_;
 wire _13814_;
 wire _13815_;
 wire _13816_;
 wire _13817_;
 wire _13818_;
 wire _13819_;
 wire _13820_;
 wire _13821_;
 wire _13822_;
 wire _13823_;
 wire _13824_;
 wire _13825_;
 wire _13826_;
 wire _13827_;
 wire _13828_;
 wire _13829_;
 wire _13830_;
 wire _13831_;
 wire _13832_;
 wire _13833_;
 wire _13834_;
 wire _13835_;
 wire _13836_;
 wire _13837_;
 wire _13838_;
 wire _13839_;
 wire _13840_;
 wire net1115;
 wire _13842_;
 wire _13843_;
 wire _13844_;
 wire _13845_;
 wire _13846_;
 wire _13847_;
 wire _13848_;
 wire _13849_;
 wire _13850_;
 wire _13851_;
 wire _13852_;
 wire _13853_;
 wire _13854_;
 wire _13855_;
 wire _13856_;
 wire _13857_;
 wire _13858_;
 wire _13859_;
 wire _13860_;
 wire _13861_;
 wire _13862_;
 wire _13863_;
 wire _13864_;
 wire _13865_;
 wire _13866_;
 wire _13867_;
 wire _13868_;
 wire _13869_;
 wire _13870_;
 wire _13871_;
 wire _13872_;
 wire _13873_;
 wire _13874_;
 wire _13875_;
 wire _13876_;
 wire _13877_;
 wire _13878_;
 wire _13879_;
 wire _13880_;
 wire _13881_;
 wire _13882_;
 wire _13883_;
 wire _13884_;
 wire _13885_;
 wire _13886_;
 wire _13887_;
 wire _13888_;
 wire _13889_;
 wire _13890_;
 wire _13891_;
 wire _13892_;
 wire _13893_;
 wire _13894_;
 wire _13895_;
 wire _13896_;
 wire _13897_;
 wire _13898_;
 wire _13899_;
 wire _13900_;
 wire _13901_;
 wire _13902_;
 wire _13903_;
 wire _13904_;
 wire _13905_;
 wire _13906_;
 wire _13907_;
 wire _13908_;
 wire _13909_;
 wire _13910_;
 wire _13911_;
 wire _13912_;
 wire _13913_;
 wire _13914_;
 wire _13915_;
 wire _13916_;
 wire _13917_;
 wire _13918_;
 wire _13919_;
 wire _13920_;
 wire _13921_;
 wire _13922_;
 wire _13923_;
 wire _13924_;
 wire _13925_;
 wire _13926_;
 wire _13927_;
 wire _13928_;
 wire _13929_;
 wire _13930_;
 wire _13931_;
 wire _13932_;
 wire _13933_;
 wire _13934_;
 wire _13935_;
 wire _13936_;
 wire _13937_;
 wire _13938_;
 wire _13939_;
 wire _13940_;
 wire _13941_;
 wire _13942_;
 wire _13943_;
 wire _13944_;
 wire _13945_;
 wire _13946_;
 wire _13947_;
 wire _13948_;
 wire _13949_;
 wire _13950_;
 wire _13951_;
 wire _13952_;
 wire _13953_;
 wire _13954_;
 wire net187;
 wire _13956_;
 wire _13957_;
 wire _13958_;
 wire _13959_;
 wire _13960_;
 wire _13961_;
 wire _13962_;
 wire _13963_;
 wire _13964_;
 wire _13965_;
 wire _13966_;
 wire _13967_;
 wire _13968_;
 wire _13969_;
 wire _13970_;
 wire _13971_;
 wire _13972_;
 wire _13973_;
 wire _13974_;
 wire _13975_;
 wire _13976_;
 wire _13977_;
 wire _13978_;
 wire net149;
 wire _13980_;
 wire _13981_;
 wire _13982_;
 wire _13983_;
 wire _13984_;
 wire _13985_;
 wire _13986_;
 wire _13987_;
 wire _13988_;
 wire _13989_;
 wire _13990_;
 wire _13991_;
 wire _13992_;
 wire _13993_;
 wire _13994_;
 wire _13995_;
 wire _13996_;
 wire _13997_;
 wire _13998_;
 wire _13999_;
 wire _14000_;
 wire _14001_;
 wire _14002_;
 wire _14003_;
 wire _14004_;
 wire _14005_;
 wire _14006_;
 wire _14007_;
 wire _14008_;
 wire _14009_;
 wire _14010_;
 wire _14011_;
 wire _14012_;
 wire _14013_;
 wire _14014_;
 wire _14015_;
 wire _14016_;
 wire _14017_;
 wire _14018_;
 wire _14019_;
 wire _14020_;
 wire _14021_;
 wire _14022_;
 wire _14023_;
 wire _14024_;
 wire _14025_;
 wire _14026_;
 wire _14027_;
 wire _14028_;
 wire _14029_;
 wire _14030_;
 wire _14031_;
 wire _14032_;
 wire _14033_;
 wire _14034_;
 wire _14035_;
 wire _14036_;
 wire _14037_;
 wire _14038_;
 wire _14039_;
 wire _14040_;
 wire _14041_;
 wire _14042_;
 wire _14043_;
 wire _14044_;
 wire _14045_;
 wire _14046_;
 wire _14047_;
 wire _14048_;
 wire _14049_;
 wire _14050_;
 wire _14051_;
 wire _14052_;
 wire _14053_;
 wire _14054_;
 wire _14055_;
 wire _14056_;
 wire _14057_;
 wire _14058_;
 wire _14059_;
 wire _14060_;
 wire _14061_;
 wire _14062_;
 wire _14063_;
 wire _14064_;
 wire _14065_;
 wire _14066_;
 wire _14067_;
 wire _14068_;
 wire _14069_;
 wire _14070_;
 wire _14071_;
 wire _14072_;
 wire _14073_;
 wire _14074_;
 wire _14075_;
 wire _14076_;
 wire _14077_;
 wire _14078_;
 wire _14079_;
 wire _14080_;
 wire _14081_;
 wire _14082_;
 wire _14083_;
 wire _14084_;
 wire _14085_;
 wire _14086_;
 wire _14087_;
 wire _14088_;
 wire _14089_;
 wire _14090_;
 wire _14091_;
 wire _14092_;
 wire _14093_;
 wire _14094_;
 wire _14095_;
 wire _14096_;
 wire _14097_;
 wire _14098_;
 wire _14099_;
 wire _14100_;
 wire _14101_;
 wire _14102_;
 wire _14103_;
 wire _14104_;
 wire _14105_;
 wire _14106_;
 wire _14107_;
 wire _14108_;
 wire _14109_;
 wire _14110_;
 wire _14111_;
 wire _14112_;
 wire _14113_;
 wire _14114_;
 wire _14115_;
 wire _14116_;
 wire _14117_;
 wire _14118_;
 wire _14119_;
 wire _14120_;
 wire _14121_;
 wire _14122_;
 wire _14123_;
 wire _14124_;
 wire _14125_;
 wire _14126_;
 wire _14127_;
 wire _14128_;
 wire _14129_;
 wire _14130_;
 wire _14131_;
 wire _14132_;
 wire _14133_;
 wire _14134_;
 wire _14135_;
 wire _14136_;
 wire _14137_;
 wire _14138_;
 wire _14139_;
 wire _14140_;
 wire _14141_;
 wire _14142_;
 wire _14143_;
 wire _14144_;
 wire _14145_;
 wire _14146_;
 wire _14147_;
 wire _14148_;
 wire _14149_;
 wire _14150_;
 wire _14151_;
 wire _14152_;
 wire _14153_;
 wire _14154_;
 wire _14155_;
 wire _14156_;
 wire _14157_;
 wire _14158_;
 wire _14159_;
 wire _14160_;
 wire _14161_;
 wire _14162_;
 wire _14163_;
 wire _14164_;
 wire _14165_;
 wire _14166_;
 wire _14167_;
 wire _14168_;
 wire _14169_;
 wire _14170_;
 wire _14171_;
 wire _14172_;
 wire _14173_;
 wire _14174_;
 wire _14175_;
 wire _14176_;
 wire _14177_;
 wire _14178_;
 wire _14179_;
 wire _14180_;
 wire _14181_;
 wire _14182_;
 wire _14183_;
 wire _14184_;
 wire _14185_;
 wire _14186_;
 wire _14187_;
 wire _14188_;
 wire _14189_;
 wire _14190_;
 wire _14191_;
 wire _14192_;
 wire _14193_;
 wire _14194_;
 wire _14195_;
 wire _14196_;
 wire _14197_;
 wire _14198_;
 wire _14199_;
 wire _14200_;
 wire _14201_;
 wire _14202_;
 wire _14203_;
 wire _14204_;
 wire _14205_;
 wire _14206_;
 wire _14207_;
 wire _14208_;
 wire _14209_;
 wire _14210_;
 wire _14211_;
 wire _14212_;
 wire _14213_;
 wire _14214_;
 wire _14215_;
 wire _14216_;
 wire _14217_;
 wire _14218_;
 wire _14219_;
 wire _14220_;
 wire _14221_;
 wire _14222_;
 wire _14223_;
 wire _14224_;
 wire _14225_;
 wire _14226_;
 wire _14227_;
 wire _14228_;
 wire _14229_;
 wire _14230_;
 wire _14231_;
 wire _14232_;
 wire _14233_;
 wire _14234_;
 wire _14235_;
 wire _14236_;
 wire _14237_;
 wire _14238_;
 wire _14239_;
 wire _14240_;
 wire _14241_;
 wire _14242_;
 wire _14243_;
 wire _14244_;
 wire _14245_;
 wire _14246_;
 wire _14247_;
 wire _14248_;
 wire _14249_;
 wire _14250_;
 wire _14251_;
 wire _14252_;
 wire _14253_;
 wire _14254_;
 wire _14255_;
 wire _14256_;
 wire _14257_;
 wire _14258_;
 wire _14259_;
 wire _14260_;
 wire _14261_;
 wire _14262_;
 wire _14263_;
 wire _14264_;
 wire _14265_;
 wire _14266_;
 wire _14267_;
 wire _14268_;
 wire _14269_;
 wire _14270_;
 wire _14271_;
 wire _14272_;
 wire _14273_;
 wire _14274_;
 wire _14275_;
 wire _14276_;
 wire _14277_;
 wire _14278_;
 wire _14279_;
 wire _14280_;
 wire _14281_;
 wire _14282_;
 wire _14283_;
 wire _14284_;
 wire _14285_;
 wire _14286_;
 wire _14287_;
 wire _14288_;
 wire _14289_;
 wire _14290_;
 wire _14291_;
 wire _14292_;
 wire _14293_;
 wire _14294_;
 wire _14295_;
 wire _14296_;
 wire _14297_;
 wire _14298_;
 wire _14299_;
 wire _14300_;
 wire _14301_;
 wire _14302_;
 wire _14303_;
 wire _14304_;
 wire _14305_;
 wire _14306_;
 wire _14307_;
 wire _14308_;
 wire _14309_;
 wire _14310_;
 wire _14311_;
 wire _14312_;
 wire _14313_;
 wire _14314_;
 wire _14315_;
 wire _14316_;
 wire _14317_;
 wire _14318_;
 wire _14319_;
 wire _14320_;
 wire _14321_;
 wire _14322_;
 wire _14323_;
 wire _14324_;
 wire _14325_;
 wire _14326_;
 wire _14327_;
 wire _14328_;
 wire _14329_;
 wire _14330_;
 wire _14331_;
 wire _14332_;
 wire _14333_;
 wire _14334_;
 wire _14335_;
 wire _14336_;
 wire _14337_;
 wire _14338_;
 wire _14339_;
 wire _14340_;
 wire _14341_;
 wire _14342_;
 wire _14343_;
 wire _14344_;
 wire _14345_;
 wire _14346_;
 wire _14347_;
 wire _14348_;
 wire _14349_;
 wire _14350_;
 wire _14351_;
 wire _14352_;
 wire _14353_;
 wire _14354_;
 wire _14355_;
 wire _14356_;
 wire _14357_;
 wire _14358_;
 wire _14359_;
 wire _14360_;
 wire _14361_;
 wire _14362_;
 wire _14363_;
 wire _14364_;
 wire _14365_;
 wire _14366_;
 wire _14367_;
 wire _14368_;
 wire _14369_;
 wire _14370_;
 wire _14371_;
 wire _14372_;
 wire _14373_;
 wire _14374_;
 wire _14375_;
 wire _14376_;
 wire _14377_;
 wire _14378_;
 wire _14379_;
 wire _14380_;
 wire _14381_;
 wire _14382_;
 wire _14383_;
 wire _14384_;
 wire _14385_;
 wire _14386_;
 wire _14387_;
 wire _14388_;
 wire _14389_;
 wire _14390_;
 wire _14391_;
 wire _14392_;
 wire _14393_;
 wire _14394_;
 wire _14395_;
 wire _14396_;
 wire _14397_;
 wire _14398_;
 wire _14399_;
 wire _14400_;
 wire _14401_;
 wire _14402_;
 wire _14403_;
 wire _14404_;
 wire _14405_;
 wire _14406_;
 wire _14407_;
 wire _14408_;
 wire _14409_;
 wire _14410_;
 wire _14411_;
 wire _14412_;
 wire _14413_;
 wire _14414_;
 wire _14415_;
 wire _14416_;
 wire _14417_;
 wire _14418_;
 wire _14419_;
 wire _14420_;
 wire _14421_;
 wire _14422_;
 wire _14423_;
 wire _14424_;
 wire _14425_;
 wire _14426_;
 wire _14427_;
 wire _14428_;
 wire _14429_;
 wire _14430_;
 wire _14431_;
 wire _14432_;
 wire _14433_;
 wire _14434_;
 wire _14435_;
 wire _14436_;
 wire _14437_;
 wire _14438_;
 wire _14439_;
 wire _14440_;
 wire _14441_;
 wire _14442_;
 wire _14443_;
 wire _14444_;
 wire _14445_;
 wire _14446_;
 wire _14447_;
 wire _14448_;
 wire _14449_;
 wire _14450_;
 wire _14451_;
 wire _14452_;
 wire _14453_;
 wire _14454_;
 wire _14455_;
 wire _14456_;
 wire _14457_;
 wire _14458_;
 wire _14459_;
 wire _14460_;
 wire _14461_;
 wire _14462_;
 wire _14463_;
 wire _14464_;
 wire _14465_;
 wire _14466_;
 wire _14467_;
 wire _14468_;
 wire _14469_;
 wire _14470_;
 wire _14471_;
 wire _14472_;
 wire _14473_;
 wire _14474_;
 wire _14475_;
 wire _14476_;
 wire _14477_;
 wire _14478_;
 wire _14479_;
 wire _14480_;
 wire _14481_;
 wire _14482_;
 wire _14483_;
 wire _14484_;
 wire _14485_;
 wire _14486_;
 wire _14487_;
 wire _14488_;
 wire _14489_;
 wire _14490_;
 wire _14491_;
 wire _14492_;
 wire _14493_;
 wire _14494_;
 wire _14495_;
 wire _14496_;
 wire _14497_;
 wire _14498_;
 wire _14499_;
 wire _14500_;
 wire _14501_;
 wire _14502_;
 wire _14503_;
 wire _14504_;
 wire _14505_;
 wire _14506_;
 wire _14507_;
 wire _14508_;
 wire _14509_;
 wire _14510_;
 wire _14511_;
 wire _14512_;
 wire _14513_;
 wire _14514_;
 wire _14515_;
 wire _14516_;
 wire _14517_;
 wire _14518_;
 wire _14519_;
 wire _14520_;
 wire _14521_;
 wire _14522_;
 wire _14523_;
 wire _14524_;
 wire _14525_;
 wire _14526_;
 wire _14527_;
 wire _14528_;
 wire _14529_;
 wire _14530_;
 wire _14531_;
 wire _14532_;
 wire _14533_;
 wire _14534_;
 wire _14535_;
 wire _14536_;
 wire _14537_;
 wire _14538_;
 wire _14539_;
 wire _14540_;
 wire _14541_;
 wire _14542_;
 wire _14543_;
 wire _14544_;
 wire _14545_;
 wire _14546_;
 wire _14547_;
 wire _14548_;
 wire _14549_;
 wire _14550_;
 wire _14551_;
 wire _14552_;
 wire _14553_;
 wire _14554_;
 wire _14555_;
 wire _14556_;
 wire _14557_;
 wire _14558_;
 wire _14559_;
 wire _14560_;
 wire _14561_;
 wire _14562_;
 wire _14563_;
 wire _14564_;
 wire _14565_;
 wire _14566_;
 wire _14567_;
 wire _14568_;
 wire _14569_;
 wire _14570_;
 wire _14571_;
 wire _14572_;
 wire _14573_;
 wire _14574_;
 wire _14575_;
 wire _14576_;
 wire _14577_;
 wire _14578_;
 wire _14579_;
 wire _14580_;
 wire _14581_;
 wire _14582_;
 wire _14583_;
 wire _14584_;
 wire _14585_;
 wire _14586_;
 wire _14587_;
 wire _14588_;
 wire _14589_;
 wire _14590_;
 wire _14591_;
 wire _14592_;
 wire _14593_;
 wire _14594_;
 wire _14595_;
 wire _14596_;
 wire _14597_;
 wire _14598_;
 wire _14599_;
 wire _14600_;
 wire _14601_;
 wire _14602_;
 wire _14603_;
 wire _14604_;
 wire _14605_;
 wire _14606_;
 wire _14607_;
 wire _14608_;
 wire _14609_;
 wire _14610_;
 wire _14611_;
 wire _14612_;
 wire _14613_;
 wire _14614_;
 wire _14615_;
 wire _14616_;
 wire _14617_;
 wire _14618_;
 wire _14619_;
 wire _14620_;
 wire _14621_;
 wire _14622_;
 wire _14623_;
 wire _14624_;
 wire _14625_;
 wire _14626_;
 wire _14627_;
 wire _14628_;
 wire _14629_;
 wire _14630_;
 wire _14631_;
 wire _14632_;
 wire _14633_;
 wire _14634_;
 wire _14635_;
 wire _14636_;
 wire _14637_;
 wire _14638_;
 wire _14639_;
 wire _14640_;
 wire _14641_;
 wire _14642_;
 wire _14643_;
 wire _14644_;
 wire _14645_;
 wire _14646_;
 wire _14647_;
 wire _14648_;
 wire _14649_;
 wire _14650_;
 wire _14651_;
 wire _14652_;
 wire _14653_;
 wire _14654_;
 wire _14655_;
 wire _14656_;
 wire _14657_;
 wire net878;
 wire _14659_;
 wire _14660_;
 wire _14661_;
 wire _14662_;
 wire _14663_;
 wire _14664_;
 wire _14665_;
 wire _14666_;
 wire _14667_;
 wire _14668_;
 wire _14669_;
 wire _14670_;
 wire _14671_;
 wire _14672_;
 wire _14673_;
 wire _14674_;
 wire _14675_;
 wire _14676_;
 wire _14677_;
 wire _14678_;
 wire _14679_;
 wire _14680_;
 wire _14681_;
 wire _14682_;
 wire _14683_;
 wire _14684_;
 wire _14685_;
 wire _14686_;
 wire _14687_;
 wire _14688_;
 wire _14689_;
 wire _14690_;
 wire _14691_;
 wire _14692_;
 wire _14693_;
 wire _14694_;
 wire _14695_;
 wire _14696_;
 wire _14697_;
 wire _14698_;
 wire _14699_;
 wire _14700_;
 wire _14701_;
 wire _14702_;
 wire _14703_;
 wire _14704_;
 wire _14705_;
 wire _14706_;
 wire _14707_;
 wire _14708_;
 wire _14709_;
 wire _14710_;
 wire _14711_;
 wire _14712_;
 wire _14713_;
 wire _14714_;
 wire _14715_;
 wire _14716_;
 wire _14717_;
 wire _14718_;
 wire _14719_;
 wire _14720_;
 wire _14721_;
 wire _14722_;
 wire _14723_;
 wire _14724_;
 wire _14725_;
 wire _14726_;
 wire net1032;
 wire _14728_;
 wire _14729_;
 wire _14730_;
 wire _14731_;
 wire _14732_;
 wire _14733_;
 wire _14734_;
 wire _14735_;
 wire _14736_;
 wire _14737_;
 wire _14738_;
 wire _14739_;
 wire _14740_;
 wire _14741_;
 wire _14742_;
 wire _14743_;
 wire _14744_;
 wire _14745_;
 wire _14746_;
 wire _14747_;
 wire _14748_;
 wire _14749_;
 wire _14750_;
 wire _14751_;
 wire _14752_;
 wire _14753_;
 wire _14754_;
 wire _14755_;
 wire _14756_;
 wire _14757_;
 wire _14758_;
 wire _14759_;
 wire _14760_;
 wire _14761_;
 wire _14762_;
 wire _14763_;
 wire _14764_;
 wire _14765_;
 wire _14766_;
 wire _14767_;
 wire _14768_;
 wire _14769_;
 wire _14770_;
 wire _14771_;
 wire _14772_;
 wire _14773_;
 wire _14774_;
 wire _14775_;
 wire _14776_;
 wire _14777_;
 wire _14778_;
 wire _14779_;
 wire _14780_;
 wire _14781_;
 wire _14782_;
 wire _14783_;
 wire _14784_;
 wire _14785_;
 wire _14786_;
 wire _14787_;
 wire _14788_;
 wire _14789_;
 wire _14790_;
 wire _14791_;
 wire _14792_;
 wire _14793_;
 wire _14794_;
 wire _14795_;
 wire _14796_;
 wire _14797_;
 wire _14798_;
 wire _14799_;
 wire _14800_;
 wire _14801_;
 wire _14802_;
 wire _14803_;
 wire _14804_;
 wire _14805_;
 wire _14806_;
 wire _14807_;
 wire _14808_;
 wire _14809_;
 wire _14810_;
 wire _14811_;
 wire _14812_;
 wire _14813_;
 wire _14814_;
 wire _14815_;
 wire _14816_;
 wire _14817_;
 wire _14818_;
 wire _14819_;
 wire _14820_;
 wire _14821_;
 wire _14822_;
 wire _14823_;
 wire _14824_;
 wire _14825_;
 wire _14826_;
 wire net883;
 wire _14828_;
 wire _14829_;
 wire _14830_;
 wire _14831_;
 wire _14832_;
 wire _14833_;
 wire _14834_;
 wire _14835_;
 wire _14836_;
 wire _14837_;
 wire _14838_;
 wire _14839_;
 wire _14840_;
 wire _14841_;
 wire _14842_;
 wire _14843_;
 wire _14844_;
 wire _14845_;
 wire _14846_;
 wire _14847_;
 wire _14848_;
 wire _14849_;
 wire _14850_;
 wire _14851_;
 wire _14852_;
 wire _14853_;
 wire _14854_;
 wire _14855_;
 wire _14856_;
 wire _14857_;
 wire _14858_;
 wire _14859_;
 wire _14860_;
 wire _14861_;
 wire _14862_;
 wire _14863_;
 wire _14864_;
 wire _14865_;
 wire _14866_;
 wire _14867_;
 wire _14868_;
 wire _14869_;
 wire _14870_;
 wire _14871_;
 wire _14872_;
 wire _14873_;
 wire _14874_;
 wire _14875_;
 wire _14876_;
 wire _14877_;
 wire _14878_;
 wire _14879_;
 wire _14880_;
 wire _14881_;
 wire _14882_;
 wire _14883_;
 wire _14884_;
 wire _14885_;
 wire _14886_;
 wire _14887_;
 wire _14888_;
 wire _14889_;
 wire _14890_;
 wire _14891_;
 wire _14892_;
 wire _14893_;
 wire _14894_;
 wire _14895_;
 wire _14896_;
 wire _14897_;
 wire _14898_;
 wire _14899_;
 wire _14900_;
 wire _14901_;
 wire _14902_;
 wire _14903_;
 wire _14904_;
 wire _14905_;
 wire _14906_;
 wire _14907_;
 wire _14908_;
 wire _14909_;
 wire _14910_;
 wire _14911_;
 wire _14912_;
 wire _14913_;
 wire _14914_;
 wire _14915_;
 wire _14916_;
 wire _14917_;
 wire _14918_;
 wire _14919_;
 wire _14920_;
 wire _14921_;
 wire _14922_;
 wire net715;
 wire _14924_;
 wire _14925_;
 wire _14926_;
 wire _14927_;
 wire _14928_;
 wire _14929_;
 wire _14930_;
 wire _14931_;
 wire _14932_;
 wire _14933_;
 wire _14934_;
 wire _14935_;
 wire _14936_;
 wire _14937_;
 wire _14938_;
 wire _14939_;
 wire _14940_;
 wire _14941_;
 wire _14942_;
 wire _14943_;
 wire _14944_;
 wire _14945_;
 wire _14946_;
 wire _14947_;
 wire _14948_;
 wire _14949_;
 wire _14950_;
 wire _14951_;
 wire _14952_;
 wire _14953_;
 wire _14954_;
 wire _14955_;
 wire _14956_;
 wire _14957_;
 wire _14958_;
 wire _14959_;
 wire _14960_;
 wire _14961_;
 wire _14962_;
 wire _14963_;
 wire _14964_;
 wire _14965_;
 wire _14966_;
 wire _14967_;
 wire _14968_;
 wire _14969_;
 wire _14970_;
 wire _14971_;
 wire _14972_;
 wire _14973_;
 wire _14974_;
 wire _14975_;
 wire _14976_;
 wire _14977_;
 wire _14978_;
 wire _14979_;
 wire _14980_;
 wire _14981_;
 wire _14982_;
 wire _14983_;
 wire _14984_;
 wire _14985_;
 wire _14986_;
 wire _14987_;
 wire _14988_;
 wire _14989_;
 wire _14990_;
 wire _14991_;
 wire _14992_;
 wire _14993_;
 wire _14994_;
 wire _14995_;
 wire _14996_;
 wire _14997_;
 wire _14998_;
 wire _14999_;
 wire _15000_;
 wire _15001_;
 wire _15002_;
 wire _15003_;
 wire _15004_;
 wire _15005_;
 wire _15006_;
 wire _15007_;
 wire _15008_;
 wire _15009_;
 wire _15010_;
 wire _15011_;
 wire _15012_;
 wire _15013_;
 wire _15014_;
 wire _15015_;
 wire _15016_;
 wire _15017_;
 wire _15018_;
 wire _15019_;
 wire _15020_;
 wire _15021_;
 wire _15022_;
 wire _15023_;
 wire _15024_;
 wire _15025_;
 wire _15026_;
 wire _15027_;
 wire _15028_;
 wire _15029_;
 wire _15030_;
 wire _15031_;
 wire _15032_;
 wire _15033_;
 wire _15034_;
 wire _15035_;
 wire _15036_;
 wire _15037_;
 wire _15038_;
 wire _15039_;
 wire _15040_;
 wire _15041_;
 wire _15042_;
 wire _15043_;
 wire _15044_;
 wire _15045_;
 wire _15046_;
 wire _15047_;
 wire _15048_;
 wire _15049_;
 wire _15050_;
 wire net843;
 wire _15052_;
 wire _15053_;
 wire _15054_;
 wire _15055_;
 wire net945;
 wire _15057_;
 wire _15058_;
 wire _15059_;
 wire _15060_;
 wire _15061_;
 wire _15062_;
 wire _15063_;
 wire _15064_;
 wire _15065_;
 wire _15066_;
 wire _15067_;
 wire _15068_;
 wire _15069_;
 wire _15070_;
 wire _15071_;
 wire _15072_;
 wire _15073_;
 wire _15074_;
 wire _15075_;
 wire _15076_;
 wire _15077_;
 wire _15078_;
 wire _15079_;
 wire _15080_;
 wire _15081_;
 wire _15082_;
 wire _15083_;
 wire _15084_;
 wire _15085_;
 wire _15086_;
 wire _15087_;
 wire _15088_;
 wire _15089_;
 wire _15090_;
 wire _15091_;
 wire _15092_;
 wire _15093_;
 wire _15094_;
 wire _15095_;
 wire _15096_;
 wire _15097_;
 wire _15098_;
 wire _15099_;
 wire _15100_;
 wire _15101_;
 wire _15102_;
 wire _15103_;
 wire _15104_;
 wire _15105_;
 wire _15106_;
 wire _15107_;
 wire _15108_;
 wire _15109_;
 wire _15110_;
 wire _15111_;
 wire _15112_;
 wire _15113_;
 wire _15114_;
 wire _15115_;
 wire _15116_;
 wire _15117_;
 wire _15118_;
 wire _15119_;
 wire _15120_;
 wire _15121_;
 wire _15122_;
 wire net599;
 wire _15124_;
 wire _15125_;
 wire _15126_;
 wire _15127_;
 wire net801;
 wire _15129_;
 wire _15130_;
 wire _15131_;
 wire _15132_;
 wire _15133_;
 wire _15134_;
 wire _15135_;
 wire _15136_;
 wire _15137_;
 wire _15138_;
 wire _15139_;
 wire _15140_;
 wire _15141_;
 wire _15142_;
 wire _15143_;
 wire _15144_;
 wire _15145_;
 wire _15146_;
 wire _15147_;
 wire _15148_;
 wire _15149_;
 wire _15150_;
 wire _15151_;
 wire _15152_;
 wire _15153_;
 wire _15154_;
 wire _15155_;
 wire _15156_;
 wire _15157_;
 wire _15158_;
 wire _15159_;
 wire _15160_;
 wire _15161_;
 wire _15162_;
 wire _15163_;
 wire _15164_;
 wire _15165_;
 wire _15166_;
 wire _15167_;
 wire _15168_;
 wire _15169_;
 wire _15170_;
 wire _15171_;
 wire _15172_;
 wire _15173_;
 wire _15174_;
 wire _15175_;
 wire _15176_;
 wire _15177_;
 wire _15178_;
 wire _15179_;
 wire _15180_;
 wire _15181_;
 wire _15182_;
 wire _15183_;
 wire _15184_;
 wire _15185_;
 wire _15186_;
 wire _15187_;
 wire _15188_;
 wire _15189_;
 wire _15190_;
 wire _15191_;
 wire _15192_;
 wire _15193_;
 wire _15194_;
 wire _15195_;
 wire _15196_;
 wire _15197_;
 wire _15198_;
 wire _15199_;
 wire net849;
 wire _15201_;
 wire _15202_;
 wire _15203_;
 wire _15204_;
 wire _15205_;
 wire _15206_;
 wire _15207_;
 wire _15208_;
 wire _15209_;
 wire _15210_;
 wire _15211_;
 wire _15212_;
 wire _15213_;
 wire _15214_;
 wire _15215_;
 wire _15216_;
 wire _15217_;
 wire _15218_;
 wire _15219_;
 wire _15220_;
 wire _15221_;
 wire _15222_;
 wire _15223_;
 wire _15224_;
 wire _15225_;
 wire _15226_;
 wire net1161;
 wire _15228_;
 wire _15229_;
 wire _15230_;
 wire _15231_;
 wire _15232_;
 wire _15233_;
 wire _15234_;
 wire _15235_;
 wire _15236_;
 wire _15237_;
 wire _15238_;
 wire _15239_;
 wire _15240_;
 wire _15241_;
 wire _15242_;
 wire _15243_;
 wire _15244_;
 wire _15245_;
 wire _15246_;
 wire _15247_;
 wire _15248_;
 wire _15249_;
 wire _15250_;
 wire _15251_;
 wire _15252_;
 wire _15253_;
 wire _15254_;
 wire _15255_;
 wire _15256_;
 wire _15257_;
 wire _15258_;
 wire _15259_;
 wire _15260_;
 wire _15261_;
 wire _15262_;
 wire _15263_;
 wire _15264_;
 wire _15265_;
 wire _15266_;
 wire _15267_;
 wire _15268_;
 wire _15269_;
 wire _15270_;
 wire _15271_;
 wire _15272_;
 wire _15273_;
 wire _15274_;
 wire _15275_;
 wire _15276_;
 wire _15277_;
 wire _15278_;
 wire _15279_;
 wire _15280_;
 wire _15281_;
 wire _15282_;
 wire _15283_;
 wire _15284_;
 wire _15285_;
 wire _15286_;
 wire _15287_;
 wire _15288_;
 wire _15289_;
 wire _15290_;
 wire _15291_;
 wire _15292_;
 wire _15293_;
 wire _15294_;
 wire _15295_;
 wire _15296_;
 wire _15297_;
 wire _15298_;
 wire _15299_;
 wire _15300_;
 wire _15301_;
 wire _15302_;
 wire _15303_;
 wire _15304_;
 wire _15305_;
 wire _15306_;
 wire _15307_;
 wire _15308_;
 wire _15309_;
 wire _15310_;
 wire _15311_;
 wire _15312_;
 wire _15313_;
 wire _15314_;
 wire _15315_;
 wire _15316_;
 wire _15317_;
 wire _15318_;
 wire _15319_;
 wire _15320_;
 wire _15321_;
 wire _15322_;
 wire _15323_;
 wire _15324_;
 wire _15325_;
 wire _15326_;
 wire _15327_;
 wire _15328_;
 wire _15329_;
 wire _15330_;
 wire _15331_;
 wire \dcnt[0] ;
 wire \dcnt[1] ;
 wire \dcnt[2] ;
 wire \dcnt[3] ;
 wire net356;
 wire ld_r;
 wire \sa00_sr[0] ;
 wire \sa00_sr[1] ;
 wire \sa00_sr[2] ;
 wire \sa00_sr[3] ;
 wire \sa00_sr[4] ;
 wire \sa00_sr[5] ;
 wire \sa00_sr[6] ;
 wire \sa00_sr[7] ;
 wire \sa01_sr[0] ;
 wire \sa01_sr[1] ;
 wire \sa01_sr[2] ;
 wire \sa01_sr[3] ;
 wire \sa01_sr[4] ;
 wire \sa01_sr[5] ;
 wire \sa01_sr[6] ;
 wire \sa01_sr[7] ;
 wire \sa02_sr[0] ;
 wire \sa02_sr[1] ;
 wire \sa02_sr[2] ;
 wire \sa02_sr[3] ;
 wire \sa02_sr[4] ;
 wire \sa02_sr[5] ;
 wire \sa02_sr[6] ;
 wire \sa02_sr[7] ;
 wire \sa03_sr[0] ;
 wire \sa03_sr[1] ;
 wire \sa03_sr[2] ;
 wire \sa03_sr[3] ;
 wire \sa03_sr[4] ;
 wire \sa03_sr[5] ;
 wire \sa03_sr[6] ;
 wire \sa03_sr[7] ;
 wire \sa10_sr[0] ;
 wire \sa10_sr[1] ;
 wire \sa10_sr[2] ;
 wire \sa10_sr[3] ;
 wire \sa10_sr[4] ;
 wire \sa10_sr[5] ;
 wire \sa10_sr[6] ;
 wire \sa10_sr[7] ;
 wire \sa10_sub[0] ;
 wire \sa10_sub[1] ;
 wire \sa10_sub[2] ;
 wire \sa10_sub[3] ;
 wire \sa10_sub[4] ;
 wire \sa10_sub[5] ;
 wire \sa10_sub[6] ;
 wire \sa10_sub[7] ;
 wire \sa11_sr[0] ;
 wire \sa11_sr[1] ;
 wire \sa11_sr[2] ;
 wire \sa11_sr[3] ;
 wire \sa11_sr[4] ;
 wire \sa11_sr[5] ;
 wire \sa11_sr[6] ;
 wire \sa11_sr[7] ;
 wire \sa12_sr[0] ;
 wire \sa12_sr[1] ;
 wire \sa12_sr[2] ;
 wire \sa12_sr[3] ;
 wire \sa12_sr[4] ;
 wire \sa12_sr[5] ;
 wire \sa12_sr[6] ;
 wire \sa12_sr[7] ;
 wire \sa20_sr[0] ;
 wire \sa20_sr[1] ;
 wire \sa20_sr[2] ;
 wire \sa20_sr[3] ;
 wire \sa20_sr[4] ;
 wire \sa20_sr[5] ;
 wire \sa20_sr[6] ;
 wire \sa20_sr[7] ;
 wire \sa20_sub[0] ;
 wire \sa20_sub[1] ;
 wire \sa20_sub[2] ;
 wire \sa20_sub[3] ;
 wire \sa20_sub[4] ;
 wire \sa20_sub[5] ;
 wire \sa20_sub[6] ;
 wire \sa20_sub[7] ;
 wire \sa21_sr[0] ;
 wire \sa21_sr[1] ;
 wire \sa21_sr[2] ;
 wire \sa21_sr[3] ;
 wire \sa21_sr[4] ;
 wire \sa21_sr[5] ;
 wire \sa21_sr[6] ;
 wire \sa21_sr[7] ;
 wire \sa21_sub[0] ;
 wire \sa21_sub[1] ;
 wire \sa21_sub[2] ;
 wire \sa21_sub[3] ;
 wire \sa21_sub[4] ;
 wire \sa21_sub[5] ;
 wire \sa21_sub[6] ;
 wire \sa21_sub[7] ;
 wire \sa30_sr[0] ;
 wire \sa30_sr[1] ;
 wire \sa30_sr[2] ;
 wire \sa30_sr[3] ;
 wire \sa30_sr[4] ;
 wire \sa30_sr[5] ;
 wire \sa30_sr[6] ;
 wire \sa30_sr[7] ;
 wire \sa30_sub[0] ;
 wire \sa30_sub[1] ;
 wire \sa30_sub[2] ;
 wire \sa30_sub[3] ;
 wire \sa30_sub[4] ;
 wire \sa30_sub[5] ;
 wire \sa30_sub[6] ;
 wire \sa30_sub[7] ;
 wire \sa31_sub[0] ;
 wire \sa31_sub[1] ;
 wire \sa31_sub[2] ;
 wire \sa31_sub[3] ;
 wire \sa31_sub[4] ;
 wire \sa31_sub[5] ;
 wire \sa31_sub[6] ;
 wire \sa31_sub[7] ;
 wire \sa32_sub[0] ;
 wire \sa32_sub[1] ;
 wire \sa32_sub[2] ;
 wire \sa32_sub[3] ;
 wire \sa32_sub[4] ;
 wire \sa32_sub[5] ;
 wire \sa32_sub[6] ;
 wire \sa32_sub[7] ;
 wire \text_in_r[0] ;
 wire \text_in_r[100] ;
 wire \text_in_r[101] ;
 wire \text_in_r[102] ;
 wire \text_in_r[103] ;
 wire \text_in_r[104] ;
 wire \text_in_r[105] ;
 wire \text_in_r[106] ;
 wire \text_in_r[107] ;
 wire \text_in_r[108] ;
 wire \text_in_r[109] ;
 wire \text_in_r[10] ;
 wire \text_in_r[110] ;
 wire \text_in_r[111] ;
 wire \text_in_r[112] ;
 wire \text_in_r[113] ;
 wire \text_in_r[114] ;
 wire \text_in_r[115] ;
 wire \text_in_r[116] ;
 wire \text_in_r[117] ;
 wire \text_in_r[118] ;
 wire \text_in_r[119] ;
 wire \text_in_r[11] ;
 wire \text_in_r[120] ;
 wire \text_in_r[121] ;
 wire \text_in_r[122] ;
 wire \text_in_r[123] ;
 wire \text_in_r[124] ;
 wire \text_in_r[125] ;
 wire \text_in_r[126] ;
 wire \text_in_r[127] ;
 wire \text_in_r[12] ;
 wire \text_in_r[13] ;
 wire \text_in_r[14] ;
 wire \text_in_r[15] ;
 wire \text_in_r[16] ;
 wire \text_in_r[17] ;
 wire \text_in_r[18] ;
 wire \text_in_r[19] ;
 wire \text_in_r[1] ;
 wire \text_in_r[20] ;
 wire \text_in_r[21] ;
 wire \text_in_r[22] ;
 wire \text_in_r[23] ;
 wire \text_in_r[24] ;
 wire \text_in_r[25] ;
 wire \text_in_r[26] ;
 wire \text_in_r[27] ;
 wire \text_in_r[28] ;
 wire \text_in_r[29] ;
 wire \text_in_r[2] ;
 wire \text_in_r[30] ;
 wire \text_in_r[31] ;
 wire \text_in_r[32] ;
 wire \text_in_r[33] ;
 wire \text_in_r[34] ;
 wire \text_in_r[35] ;
 wire \text_in_r[36] ;
 wire \text_in_r[37] ;
 wire \text_in_r[38] ;
 wire \text_in_r[39] ;
 wire \text_in_r[3] ;
 wire \text_in_r[40] ;
 wire \text_in_r[41] ;
 wire \text_in_r[42] ;
 wire \text_in_r[43] ;
 wire \text_in_r[44] ;
 wire \text_in_r[45] ;
 wire \text_in_r[46] ;
 wire \text_in_r[47] ;
 wire \text_in_r[48] ;
 wire \text_in_r[49] ;
 wire \text_in_r[4] ;
 wire \text_in_r[50] ;
 wire \text_in_r[51] ;
 wire \text_in_r[52] ;
 wire \text_in_r[53] ;
 wire \text_in_r[54] ;
 wire \text_in_r[55] ;
 wire \text_in_r[56] ;
 wire \text_in_r[57] ;
 wire \text_in_r[58] ;
 wire \text_in_r[59] ;
 wire \text_in_r[5] ;
 wire \text_in_r[60] ;
 wire \text_in_r[61] ;
 wire \text_in_r[62] ;
 wire \text_in_r[63] ;
 wire \text_in_r[64] ;
 wire \text_in_r[65] ;
 wire \text_in_r[66] ;
 wire \text_in_r[67] ;
 wire \text_in_r[68] ;
 wire \text_in_r[69] ;
 wire \text_in_r[6] ;
 wire \text_in_r[70] ;
 wire \text_in_r[71] ;
 wire \text_in_r[72] ;
 wire \text_in_r[73] ;
 wire \text_in_r[74] ;
 wire \text_in_r[75] ;
 wire \text_in_r[76] ;
 wire \text_in_r[77] ;
 wire \text_in_r[78] ;
 wire \text_in_r[79] ;
 wire \text_in_r[7] ;
 wire \text_in_r[80] ;
 wire \text_in_r[81] ;
 wire \text_in_r[82] ;
 wire \text_in_r[83] ;
 wire \text_in_r[84] ;
 wire \text_in_r[85] ;
 wire \text_in_r[86] ;
 wire \text_in_r[87] ;
 wire \text_in_r[88] ;
 wire \text_in_r[89] ;
 wire \text_in_r[8] ;
 wire \text_in_r[90] ;
 wire \text_in_r[91] ;
 wire \text_in_r[92] ;
 wire \text_in_r[93] ;
 wire \text_in_r[94] ;
 wire \text_in_r[95] ;
 wire \text_in_r[96] ;
 wire \text_in_r[97] ;
 wire \text_in_r[98] ;
 wire \text_in_r[99] ;
 wire \text_in_r[9] ;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire \u0.r0.out[24] ;
 wire \u0.r0.out[25] ;
 wire \u0.r0.out[26] ;
 wire \u0.r0.out[27] ;
 wire \u0.r0.out[28] ;
 wire \u0.r0.out[29] ;
 wire \u0.r0.out[30] ;
 wire \u0.r0.out[31] ;
 wire \u0.r0.rcnt[0] ;
 wire \u0.r0.rcnt[1] ;
 wire \u0.r0.rcnt[2] ;
 wire \u0.r0.rcnt[3] ;
 wire \u0.r0.rcnt_next[0] ;
 wire \u0.r0.rcnt_next[1] ;
 wire \u0.subword[0] ;
 wire \u0.subword[10] ;
 wire \u0.subword[11] ;
 wire \u0.subword[12] ;
 wire \u0.subword[13] ;
 wire \u0.subword[14] ;
 wire \u0.subword[15] ;
 wire \u0.subword[16] ;
 wire \u0.subword[17] ;
 wire \u0.subword[18] ;
 wire \u0.subword[19] ;
 wire \u0.subword[1] ;
 wire \u0.subword[20] ;
 wire \u0.subword[21] ;
 wire \u0.subword[22] ;
 wire \u0.subword[23] ;
 wire \u0.subword[24] ;
 wire \u0.subword[25] ;
 wire \u0.subword[26] ;
 wire \u0.subword[27] ;
 wire \u0.subword[28] ;
 wire \u0.subword[29] ;
 wire \u0.subword[2] ;
 wire \u0.subword[30] ;
 wire \u0.subword[31] ;
 wire \u0.subword[3] ;
 wire \u0.subword[4] ;
 wire \u0.subword[5] ;
 wire \u0.subword[6] ;
 wire \u0.subword[7] ;
 wire \u0.subword[8] ;
 wire \u0.subword[9] ;
 wire \u0.tmp_w[0] ;
 wire \u0.tmp_w[10] ;
 wire \u0.tmp_w[11] ;
 wire \u0.tmp_w[12] ;
 wire \u0.tmp_w[13] ;
 wire \u0.tmp_w[14] ;
 wire \u0.tmp_w[15] ;
 wire \u0.tmp_w[16] ;
 wire \u0.tmp_w[17] ;
 wire \u0.tmp_w[18] ;
 wire \u0.tmp_w[19] ;
 wire \u0.tmp_w[1] ;
 wire \u0.tmp_w[20] ;
 wire \u0.tmp_w[21] ;
 wire \u0.tmp_w[22] ;
 wire \u0.tmp_w[23] ;
 wire \u0.tmp_w[24] ;
 wire \u0.tmp_w[25] ;
 wire \u0.tmp_w[26] ;
 wire \u0.tmp_w[27] ;
 wire \u0.tmp_w[28] ;
 wire \u0.tmp_w[29] ;
 wire \u0.tmp_w[2] ;
 wire \u0.tmp_w[30] ;
 wire \u0.tmp_w[31] ;
 wire \u0.tmp_w[3] ;
 wire \u0.tmp_w[4] ;
 wire \u0.tmp_w[5] ;
 wire \u0.tmp_w[6] ;
 wire \u0.tmp_w[7] ;
 wire \u0.tmp_w[8] ;
 wire \u0.tmp_w[9] ;
 wire \u0.w[0][0] ;
 wire \u0.w[0][10] ;
 wire \u0.w[0][11] ;
 wire \u0.w[0][12] ;
 wire \u0.w[0][13] ;
 wire \u0.w[0][14] ;
 wire \u0.w[0][15] ;
 wire \u0.w[0][16] ;
 wire \u0.w[0][17] ;
 wire \u0.w[0][18] ;
 wire \u0.w[0][19] ;
 wire \u0.w[0][1] ;
 wire \u0.w[0][20] ;
 wire \u0.w[0][21] ;
 wire \u0.w[0][22] ;
 wire \u0.w[0][23] ;
 wire \u0.w[0][24] ;
 wire \u0.w[0][25] ;
 wire \u0.w[0][26] ;
 wire \u0.w[0][27] ;
 wire \u0.w[0][28] ;
 wire \u0.w[0][29] ;
 wire \u0.w[0][2] ;
 wire \u0.w[0][30] ;
 wire \u0.w[0][31] ;
 wire \u0.w[0][3] ;
 wire \u0.w[0][4] ;
 wire \u0.w[0][5] ;
 wire \u0.w[0][6] ;
 wire \u0.w[0][7] ;
 wire \u0.w[0][8] ;
 wire \u0.w[0][9] ;
 wire \u0.w[1][0] ;
 wire \u0.w[1][10] ;
 wire \u0.w[1][11] ;
 wire \u0.w[1][12] ;
 wire \u0.w[1][13] ;
 wire \u0.w[1][14] ;
 wire \u0.w[1][15] ;
 wire \u0.w[1][16] ;
 wire \u0.w[1][17] ;
 wire \u0.w[1][18] ;
 wire \u0.w[1][19] ;
 wire \u0.w[1][1] ;
 wire \u0.w[1][20] ;
 wire \u0.w[1][21] ;
 wire \u0.w[1][22] ;
 wire \u0.w[1][23] ;
 wire \u0.w[1][24] ;
 wire \u0.w[1][25] ;
 wire \u0.w[1][26] ;
 wire \u0.w[1][27] ;
 wire \u0.w[1][28] ;
 wire \u0.w[1][29] ;
 wire \u0.w[1][2] ;
 wire \u0.w[1][30] ;
 wire \u0.w[1][31] ;
 wire \u0.w[1][3] ;
 wire \u0.w[1][4] ;
 wire \u0.w[1][5] ;
 wire \u0.w[1][6] ;
 wire \u0.w[1][7] ;
 wire \u0.w[1][8] ;
 wire \u0.w[1][9] ;
 wire \u0.w[2][0] ;
 wire \u0.w[2][10] ;
 wire \u0.w[2][11] ;
 wire \u0.w[2][12] ;
 wire \u0.w[2][13] ;
 wire \u0.w[2][14] ;
 wire \u0.w[2][15] ;
 wire \u0.w[2][16] ;
 wire \u0.w[2][17] ;
 wire \u0.w[2][18] ;
 wire \u0.w[2][19] ;
 wire \u0.w[2][1] ;
 wire \u0.w[2][20] ;
 wire \u0.w[2][21] ;
 wire \u0.w[2][22] ;
 wire \u0.w[2][23] ;
 wire \u0.w[2][24] ;
 wire \u0.w[2][25] ;
 wire \u0.w[2][26] ;
 wire \u0.w[2][27] ;
 wire \u0.w[2][28] ;
 wire \u0.w[2][29] ;
 wire \u0.w[2][2] ;
 wire \u0.w[2][30] ;
 wire \u0.w[2][31] ;
 wire \u0.w[2][3] ;
 wire \u0.w[2][4] ;
 wire \u0.w[2][5] ;
 wire \u0.w[2][6] ;
 wire \u0.w[2][7] ;
 wire \u0.w[2][8] ;
 wire \u0.w[2][9] ;
 wire net103;
 wire net105;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net123;
 wire net124;
 wire net125;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net10;
 wire net11;
 wire net17;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net30;
 wire net31;
 wire net33;
 wire net34;
 wire net35;
 wire net38;
 wire net40;
 wire net41;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net50;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net104;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net142;
 wire net147;
 wire net148;
 wire net150;
 wire net151;
 wire net158;
 wire net163;
 wire net164;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net172;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net198;
 wire net199;
 wire net201;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire clknet_leaf_0_clk;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_leaf_45_clk;
 wire clknet_leaf_46_clk;
 wire clknet_leaf_47_clk;
 wire clknet_leaf_48_clk;
 wire clknet_leaf_49_clk;
 wire clknet_leaf_50_clk;
 wire clknet_leaf_51_clk;
 wire clknet_leaf_52_clk;
 wire clknet_leaf_53_clk;
 wire clknet_leaf_54_clk;
 wire clknet_leaf_55_clk;
 wire clknet_leaf_56_clk;
 wire clknet_leaf_57_clk;
 wire clknet_leaf_58_clk;
 wire clknet_leaf_59_clk;
 wire clknet_leaf_60_clk;
 wire clknet_leaf_61_clk;
 wire clknet_leaf_62_clk;
 wire clknet_leaf_63_clk;
 wire clknet_leaf_64_clk;
 wire clknet_leaf_65_clk;
 wire clknet_leaf_66_clk;
 wire clknet_leaf_67_clk;
 wire clknet_leaf_68_clk;
 wire clknet_leaf_69_clk;
 wire clknet_leaf_70_clk;
 wire clknet_leaf_71_clk;
 wire clknet_leaf_72_clk;
 wire clknet_leaf_73_clk;
 wire clknet_leaf_74_clk;
 wire clknet_leaf_75_clk;
 wire clknet_leaf_76_clk;
 wire clknet_leaf_77_clk;
 wire clknet_leaf_78_clk;
 wire clknet_leaf_79_clk;
 wire clknet_leaf_80_clk;
 wire clknet_leaf_81_clk;
 wire clknet_leaf_82_clk;
 wire clknet_leaf_83_clk;
 wire clknet_leaf_84_clk;
 wire clknet_leaf_85_clk;
 wire clknet_leaf_86_clk;
 wire clknet_leaf_87_clk;
 wire clknet_leaf_88_clk;
 wire clknet_leaf_89_clk;
 wire clknet_leaf_90_clk;
 wire clknet_leaf_91_clk;
 wire clknet_leaf_92_clk;
 wire clknet_leaf_93_clk;
 wire clknet_leaf_94_clk;
 wire clknet_leaf_95_clk;
 wire clknet_leaf_96_clk;
 wire clknet_leaf_97_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net600;
 wire net1224;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net616;
 wire net618;
 wire net619;
 wire net620;
 wire net629;
 wire net630;
 wire net631;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net645;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net654;
 wire net655;
 wire net656;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net725;
 wire net726;
 wire net727;
 wire net734;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net783;
 wire net784;
 wire net785;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net796;
 wire net797;
 wire net798;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net825;
 wire net826;
 wire net827;
 wire net830;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net848;
 wire net871;
 wire net885;
 wire net896;
 wire net897;
 wire net898;
 wire net901;
 wire net902;
 wire net909;
 wire net910;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net931;
 wire net932;
 wire net943;
 wire net944;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net1001;
 wire net1002;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1033;
 wire net1036;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1056;
 wire net1057;
 wire net1068;
 wire net1069;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1088;
 wire net1089;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1112;
 wire net1114;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1163;
 wire net1164;
 wire net1167;
 wire net1174;
 wire net1175;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1200;
 wire net1201;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1;
 wire net615;
 wire net621;
 wire net673;
 wire net698;
 wire net705;
 wire net706;
 wire net707;
 wire net714;
 wire net718;
 wire net719;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net735;
 wire net802;
 wire net803;
 wire net805;
 wire net807;
 wire net829;
 wire net831;
 wire net832;
 wire net835;
 wire net844;
 wire net847;
 wire net850;
 wire net851;
 wire net852;
 wire net879;
 wire net911;
 wire net915;
 wire net916;
 wire net918;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net955;
 wire net956;
 wire net992;
 wire net993;
 wire net997;
 wire net999;
 wire net1000;
 wire net1003;
 wire net1004;
 wire net1030;
 wire net1037;
 wire net1038;
 wire net1045;
 wire net1046;
 wire net1084;
 wire net1085;
 wire net1116;
 wire net1124;
 wire net1144;
 wire net1147;
 wire net1159;
 wire net1165;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1182;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1197;
 wire net1198;
 wire net1202;
 wire net1203;
 wire net1209;
 wire net1226;
 wire net1227;
 wire net1230;
 wire net1234;
 wire net1235;
 wire net1240;
 wire net1241;

 BUF_X16 _15332_ (.A(net226),
    .Z(_06216_));
 INV_X8 _15333_ (.A(_06216_),
    .ZN(_06217_));
 BUF_X8 _15334_ (.A(_06217_),
    .Z(_06218_));
 NOR2_X2 _15335_ (.A1(_06218_),
    .A2(net72),
    .ZN(_06219_));
 BUF_X8 _15336_ (.A(_06217_),
    .Z(_06220_));
 CLKBUF_X3 _15337_ (.A(\u0.w[0][19] ),
    .Z(_06221_));
 BUF_X4 _15338_ (.A(\u0.w[1][19] ),
    .Z(_06222_));
 XNOR2_X2 _15339_ (.A(_06221_),
    .B(_06222_),
    .ZN(_06223_));
 AND2_X1 _15340_ (.A1(_06220_),
    .A2(_06223_),
    .ZN(_06224_));
 BUF_X8 _15341_ (.A(_06216_),
    .Z(_06225_));
 BUF_X8 _15342_ (.A(_06225_),
    .Z(_06226_));
 NOR2_X1 _15343_ (.A1(net16),
    .A2(_06223_),
    .ZN(_06227_));
 CLKBUF_X3 _15344_ (.A(\u0.w[2][19] ),
    .Z(_06228_));
 BUF_X4 _15345_ (.A(\u0.tmp_w[19] ),
    .Z(_06229_));
 XNOR2_X1 _15346_ (.A(_06229_),
    .B(\u0.subword[19] ),
    .ZN(_06230_));
 XNOR2_X1 _15347_ (.A(_06228_),
    .B(_06230_),
    .ZN(_06231_));
 MUX2_X2 _15348_ (.A(_06224_),
    .B(_06227_),
    .S(_06231_),
    .Z(_06232_));
 OR2_X2 _15349_ (.A1(_06219_),
    .A2(_06232_),
    .ZN(_06233_));
 INV_X1 _15350_ (.A(_06233_),
    .ZN(_06234_));
 BUF_X4 _15351_ (.A(_06234_),
    .Z(_06235_));
 BUF_X4 _15352_ (.A(_06235_),
    .Z(_06236_));
 BUF_X4 _15353_ (.A(_06236_),
    .Z(_06237_));
 CLKBUF_X3 _15354_ (.A(_06237_),
    .Z(_06238_));
 CLKBUF_X3 _15355_ (.A(_06238_),
    .Z(_00390_));
 BUF_X8 _15356_ (.A(_06218_),
    .Z(_06239_));
 NOR2_X2 _15357_ (.A1(_06239_),
    .A2(net69),
    .ZN(_06240_));
 BUF_X4 _15358_ (.A(\u0.w[0][16] ),
    .Z(_06241_));
 BUF_X4 _15359_ (.A(\u0.w[1][16] ),
    .Z(_06242_));
 XNOR2_X2 _15360_ (.A(_06241_),
    .B(_06242_),
    .ZN(_06243_));
 AND2_X1 _15361_ (.A1(_06218_),
    .A2(_06243_),
    .ZN(_06244_));
 BUF_X8 _15362_ (.A(_06225_),
    .Z(_06245_));
 NOR2_X1 _15363_ (.A1(_06245_),
    .A2(_06243_),
    .ZN(_06246_));
 BUF_X4 _15364_ (.A(\u0.w[2][16] ),
    .Z(_06247_));
 BUF_X1 rebuffer84 (.A(\u0.tmp_w[16] ),
    .Z(net568));
 XNOR2_X2 _15366_ (.A(\u0.tmp_w[16] ),
    .B(\u0.subword[16] ),
    .ZN(_06249_));
 XNOR2_X2 _15367_ (.A(_06249_),
    .B(_06247_),
    .ZN(_06250_));
 MUX2_X2 _15368_ (.A(_06244_),
    .B(_06246_),
    .S(_06250_),
    .Z(_06251_));
 NOR2_X4 _15369_ (.A1(_06251_),
    .A2(_06240_),
    .ZN(_06252_));
 INV_X8 _15370_ (.A(net517),
    .ZN(_06253_));
 BUF_X16 _15371_ (.A(_06253_),
    .Z(_14664_));
 NOR2_X4 _15372_ (.A1(_06239_),
    .A2(net70),
    .ZN(_06254_));
 CLKBUF_X3 _15373_ (.A(\u0.w[0][17] ),
    .Z(_06255_));
 BUF_X4 _15374_ (.A(\u0.w[1][17] ),
    .Z(_06256_));
 XNOR2_X2 _15375_ (.A(_06255_),
    .B(_06256_),
    .ZN(_06257_));
 AND2_X1 _15376_ (.A1(_06220_),
    .A2(_06257_),
    .ZN(_06258_));
 NOR2_X1 _15377_ (.A1(_06245_),
    .A2(_06257_),
    .ZN(_06259_));
 BUF_X4 _15378_ (.A(\u0.w[2][17] ),
    .Z(_06260_));
 BUF_X8 clone134 (.A(net632),
    .Z(net628));
 XNOR2_X2 _15380_ (.A(\u0.tmp_w[17] ),
    .B(\u0.subword[17] ),
    .ZN(_06262_));
 XNOR2_X2 _15381_ (.A(_06262_),
    .B(_06260_),
    .ZN(_06263_));
 MUX2_X2 _15382_ (.A(_06258_),
    .B(_06259_),
    .S(_06263_),
    .Z(_06264_));
 NOR2_X4 _15383_ (.A1(_06264_),
    .A2(_06254_),
    .ZN(_06265_));
 INV_X8 _15384_ (.A(net505),
    .ZN(_14669_));
 BUF_X8 _15385_ (.A(_06239_),
    .Z(_06266_));
 BUF_X8 _15386_ (.A(_06266_),
    .Z(_06267_));
 CLKBUF_X3 _15387_ (.A(\u0.tmp_w[21] ),
    .Z(_06268_));
 CLKBUF_X3 _15388_ (.A(\u0.w[0][21] ),
    .Z(_06269_));
 BUF_X4 _15389_ (.A(\u0.w[1][21] ),
    .Z(_06270_));
 XOR2_X2 _15390_ (.A(_06269_),
    .B(_06270_),
    .Z(_06271_));
 BUF_X4 _15391_ (.A(\u0.w[2][21] ),
    .Z(_06272_));
 XNOR2_X1 _15392_ (.A(_06272_),
    .B(\u0.subword[21] ),
    .ZN(_06273_));
 XNOR2_X1 _15393_ (.A(_06271_),
    .B(_06273_),
    .ZN(_06274_));
 XNOR2_X1 _15394_ (.A(_06268_),
    .B(_06274_),
    .ZN(_06275_));
 NAND2_X1 _15395_ (.A1(_06267_),
    .A2(_06275_),
    .ZN(_06276_));
 OAI21_X4 _15396_ (.A(_06276_),
    .B1(net75),
    .B2(_06267_),
    .ZN(_06277_));
 INV_X4 _15397_ (.A(_06277_),
    .ZN(_06278_));
 CLKBUF_X3 _15398_ (.A(_06278_),
    .Z(_00392_));
 BUF_X4 _15399_ (.A(_06245_),
    .Z(_06279_));
 AND2_X1 _15400_ (.A1(_06279_),
    .A2(net74),
    .ZN(_06280_));
 CLKBUF_X3 _15401_ (.A(\u0.w[0][20] ),
    .Z(_06281_));
 BUF_X4 _15402_ (.A(\u0.w[1][20] ),
    .Z(_06282_));
 XNOR2_X2 _15403_ (.A(_06281_),
    .B(_06282_),
    .ZN(_06283_));
 BUF_X4 _15404_ (.A(\u0.w[2][20] ),
    .Z(_06284_));
 BUF_X2 _15405_ (.A(\u0.tmp_w[20] ),
    .Z(_06285_));
 XNOR2_X1 _15406_ (.A(_06285_),
    .B(\u0.subword[20] ),
    .ZN(_06286_));
 XNOR2_X1 _15407_ (.A(_06284_),
    .B(_06286_),
    .ZN(_06287_));
 XNOR2_X2 _15408_ (.A(_06283_),
    .B(_06287_),
    .ZN(_06288_));
 AOI21_X4 _15409_ (.A(_06280_),
    .B1(_06288_),
    .B2(_06239_),
    .ZN(_06289_));
 INV_X2 _15410_ (.A(_06289_),
    .ZN(_06290_));
 BUF_X4 _15411_ (.A(_06290_),
    .Z(_06291_));
 CLKBUF_X3 _15412_ (.A(_06291_),
    .Z(_06292_));
 CLKBUF_X3 _15413_ (.A(_06292_),
    .Z(_06293_));
 CLKBUF_X3 _15414_ (.A(_06293_),
    .Z(_00391_));
 NAND2_X1 _15415_ (.A1(_06245_),
    .A2(net71),
    .ZN(_06294_));
 BUF_X4 _15416_ (.A(\u0.tmp_w[18] ),
    .Z(_06295_));
 BUF_X8 _15417_ (.A(\u0.w[0][18] ),
    .Z(_06296_));
 BUF_X4 _15418_ (.A(\u0.w[1][18] ),
    .Z(_06297_));
 XOR2_X2 _15419_ (.A(_06296_),
    .B(_06297_),
    .Z(_06298_));
 BUF_X8 _15420_ (.A(\u0.w[2][18] ),
    .Z(_06299_));
 BUF_X1 _15421_ (.A(_00408_),
    .Z(_06300_));
 NOR2_X1 _15422_ (.A1(_06299_),
    .A2(_06300_),
    .ZN(_06301_));
 NAND4_X1 _15423_ (.A1(_06217_),
    .A2(_06295_),
    .A3(_06298_),
    .A4(_06301_),
    .ZN(_06302_));
 INV_X1 _15424_ (.A(_06300_),
    .ZN(_06303_));
 NOR2_X1 _15425_ (.A1(_06216_),
    .A2(_06295_),
    .ZN(_06304_));
 NAND4_X1 _15426_ (.A1(_06299_),
    .A2(_06303_),
    .A3(_06298_),
    .A4(_06304_),
    .ZN(_06305_));
 INV_X2 _15427_ (.A(_06299_),
    .ZN(_06306_));
 NAND4_X1 _15428_ (.A1(_06306_),
    .A2(_06300_),
    .A3(_06298_),
    .A4(_06304_),
    .ZN(_06307_));
 INV_X1 _15429_ (.A(_06295_),
    .ZN(_06308_));
 XNOR2_X2 _15430_ (.A(_06297_),
    .B(_06296_),
    .ZN(_06309_));
 NAND2_X1 _15431_ (.A1(_06299_),
    .A2(_06300_),
    .ZN(_06310_));
 OR4_X4 _15432_ (.A1(_06216_),
    .A2(_06308_),
    .A3(_06309_),
    .A4(_06310_),
    .ZN(_06311_));
 AND4_X4 _15433_ (.A1(_06302_),
    .A2(_06305_),
    .A3(_06307_),
    .A4(_06311_),
    .ZN(_06312_));
 AND2_X1 _15434_ (.A1(_06301_),
    .A2(_06304_),
    .ZN(_06313_));
 NOR4_X1 _15435_ (.A1(_06225_),
    .A2(_06308_),
    .A3(_06306_),
    .A4(_06300_),
    .ZN(_06314_));
 OAI21_X1 _15436_ (.A(_06309_),
    .B1(_06313_),
    .B2(_06314_),
    .ZN(_06315_));
 NOR4_X1 _15437_ (.A1(_06225_),
    .A2(_06308_),
    .A3(_06299_),
    .A4(_06303_),
    .ZN(_06316_));
 NOR3_X1 _15438_ (.A1(_06225_),
    .A2(_06295_),
    .A3(_06310_),
    .ZN(_06317_));
 OAI21_X1 _15439_ (.A(_06309_),
    .B1(_06316_),
    .B2(_06317_),
    .ZN(_06318_));
 AND4_X4 _15440_ (.A1(_06312_),
    .A2(_06294_),
    .A3(_06315_),
    .A4(_06318_),
    .ZN(_06319_));
 BUF_X2 rebuffer736 (.A(_14925_),
    .Z(net1199));
 INV_X8 _15442_ (.A(_06319_),
    .ZN(_06321_));
 BUF_X4 _15443_ (.A(_06321_),
    .Z(_06322_));
 BUF_X8 _15444_ (.A(_06322_),
    .Z(_06323_));
 BUF_X8 _15445_ (.A(_06323_),
    .Z(_14683_));
 NOR2_X4 _15446_ (.A1(_06239_),
    .A2(net19),
    .ZN(_06324_));
 BUF_X4 _15447_ (.A(\u0.w[0][0] ),
    .Z(_06325_));
 BUF_X4 _15448_ (.A(\u0.w[1][0] ),
    .Z(_06326_));
 XNOR2_X2 _15449_ (.A(_06325_),
    .B(_06326_),
    .ZN(_06327_));
 AND2_X1 _15450_ (.A1(_06220_),
    .A2(_06327_),
    .ZN(_06328_));
 NOR2_X1 _15451_ (.A1(_06226_),
    .A2(_06327_),
    .ZN(_06329_));
 BUF_X4 _15452_ (.A(\u0.w[2][0] ),
    .Z(_06330_));
 BUF_X1 rebuffer620 (.A(_06475_),
    .Z(net1225));
 XNOR2_X2 _15454_ (.A(\u0.subword[0] ),
    .B(\u0.tmp_w[0] ),
    .ZN(_06332_));
 XNOR2_X1 _15455_ (.A(_06330_),
    .B(_06332_),
    .ZN(_06333_));
 MUX2_X2 _15456_ (.A(_06328_),
    .B(_06329_),
    .S(_06333_),
    .Z(_06334_));
 NOR2_X4 _15457_ (.A1(_06334_),
    .A2(_06324_),
    .ZN(_06335_));
 INV_X8 _15458_ (.A(net1209),
    .ZN(_06336_));
 BUF_X1 rebuffer703 (.A(_08004_),
    .Z(net1166));
 BUF_X16 _15460_ (.A(_06336_),
    .Z(_14732_));
 NOR2_X4 _15461_ (.A1(_06239_),
    .A2(net73),
    .ZN(_06338_));
 BUF_X8 _15462_ (.A(_06226_),
    .Z(_06339_));
 BUF_X4 _15463_ (.A(\u0.w[0][1] ),
    .Z(_06340_));
 BUF_X4 _15464_ (.A(\u0.w[1][1] ),
    .Z(_06341_));
 XOR2_X2 _15465_ (.A(_06340_),
    .B(_06341_),
    .Z(_06342_));
 NOR2_X1 _15466_ (.A1(_06339_),
    .A2(_06342_),
    .ZN(_06343_));
 XNOR2_X2 _15467_ (.A(_06340_),
    .B(_06341_),
    .ZN(_06344_));
 NOR2_X1 _15468_ (.A1(_06339_),
    .A2(_06344_),
    .ZN(_06345_));
 BUF_X4 _15469_ (.A(\u0.w[2][1] ),
    .Z(_06346_));
 BUF_X1 rebuffer273 (.A(\u0.subword[1] ),
    .Z(net828));
 XNOR2_X2 _15471_ (.A(\u0.subword[1] ),
    .B(\u0.tmp_w[1] ),
    .ZN(_06348_));
 XNOR2_X2 _15472_ (.A(_06346_),
    .B(_06348_),
    .ZN(_06349_));
 MUX2_X2 _15473_ (.A(_06343_),
    .B(_06345_),
    .S(_06349_),
    .Z(_06350_));
 NOR2_X4 _15474_ (.A1(_06350_),
    .A2(_06338_),
    .ZN(_06351_));
 INV_X8 _15475_ (.A(net614),
    .ZN(_06352_));
 BUF_X16 _15476_ (.A(_06352_),
    .Z(_14737_));
 NAND2_X1 _15477_ (.A1(_06245_),
    .A2(net84),
    .ZN(_06353_));
 BUF_X4 _15478_ (.A(\u0.tmp_w[2] ),
    .Z(_06354_));
 BUF_X8 _15479_ (.A(\u0.w[0][2] ),
    .Z(_06355_));
 BUF_X8 _15480_ (.A(\u0.w[1][2] ),
    .Z(_06356_));
 XOR2_X2 _15481_ (.A(_06355_),
    .B(_06356_),
    .Z(_06357_));
 BUF_X4 _15482_ (.A(\u0.w[2][2] ),
    .Z(_06358_));
 BUF_X2 _15483_ (.A(_00409_),
    .Z(_06359_));
 NOR2_X1 _15484_ (.A1(_06358_),
    .A2(_06359_),
    .ZN(_06360_));
 NAND4_X1 _15485_ (.A1(_06220_),
    .A2(_06354_),
    .A3(_06357_),
    .A4(_06360_),
    .ZN(_06361_));
 INV_X1 _15486_ (.A(_06359_),
    .ZN(_06362_));
 NOR2_X2 _15487_ (.A1(_06216_),
    .A2(_06354_),
    .ZN(_06363_));
 NAND4_X1 _15488_ (.A1(_06358_),
    .A2(_06362_),
    .A3(_06357_),
    .A4(_06363_),
    .ZN(_06364_));
 INV_X2 _15489_ (.A(_06358_),
    .ZN(_06365_));
 NAND4_X1 _15490_ (.A1(_06365_),
    .A2(_06359_),
    .A3(_06357_),
    .A4(_06363_),
    .ZN(_06366_));
 INV_X2 _15491_ (.A(_06354_),
    .ZN(_06367_));
 XNOR2_X2 _15492_ (.A(_06356_),
    .B(_06355_),
    .ZN(_06368_));
 NAND2_X1 _15493_ (.A1(\u0.w[2][2] ),
    .A2(_06359_),
    .ZN(_06369_));
 OR4_X2 _15494_ (.A1(net6),
    .A2(_06367_),
    .A3(_06368_),
    .A4(_06369_),
    .ZN(_06370_));
 AND4_X4 _15495_ (.A1(_06370_),
    .A2(_06364_),
    .A3(_06366_),
    .A4(_06361_),
    .ZN(_06371_));
 AND2_X1 _15496_ (.A1(_06360_),
    .A2(_06363_),
    .ZN(_06372_));
 NOR4_X1 _15497_ (.A1(_06226_),
    .A2(_06367_),
    .A3(_06365_),
    .A4(_06359_),
    .ZN(_06373_));
 OAI21_X1 _15498_ (.A(_06368_),
    .B1(_06372_),
    .B2(_06373_),
    .ZN(_06374_));
 NOR4_X1 _15499_ (.A1(net16),
    .A2(_06367_),
    .A3(_06358_),
    .A4(_06362_),
    .ZN(_06375_));
 NOR3_X1 _15500_ (.A1(net16),
    .A2(_06354_),
    .A3(_06369_),
    .ZN(_06376_));
 OAI21_X1 _15501_ (.A(net1162),
    .B1(_06375_),
    .B2(_06376_),
    .ZN(_06377_));
 AND4_X4 _15502_ (.A1(_06353_),
    .A2(_06371_),
    .A3(_06374_),
    .A4(_06377_),
    .ZN(_06378_));
 BUF_X8 _15503_ (.A(_06378_),
    .Z(_06379_));
 INV_X4 _15504_ (.A(_06379_),
    .ZN(_06380_));
 BUF_X8 _15505_ (.A(_06380_),
    .Z(_06381_));
 BUF_X8 _15506_ (.A(_06381_),
    .Z(_06382_));
 BUF_X4 _15507_ (.A(_06382_),
    .Z(_06383_));
 BUF_X4 _15508_ (.A(_06383_),
    .Z(_14751_));
 OR2_X1 _15509_ (.A1(_06218_),
    .A2(net116),
    .ZN(_06384_));
 BUF_X4 _15510_ (.A(_06384_),
    .Z(_06385_));
 BUF_X4 _15511_ (.A(\u0.w[0][3] ),
    .Z(_06386_));
 BUF_X4 _15512_ (.A(\u0.w[1][3] ),
    .Z(_06387_));
 XNOR2_X2 _15513_ (.A(_06386_),
    .B(_06387_),
    .ZN(_06388_));
 NAND2_X1 _15514_ (.A1(_06220_),
    .A2(_06388_),
    .ZN(_06389_));
 XOR2_X2 _15515_ (.A(_06386_),
    .B(_06387_),
    .Z(_06390_));
 NAND2_X1 _15516_ (.A1(_06220_),
    .A2(_06390_),
    .ZN(_06391_));
 BUF_X4 _15517_ (.A(\u0.w[2][3] ),
    .Z(_06392_));
 BUF_X4 _15518_ (.A(\u0.tmp_w[3] ),
    .Z(_06393_));
 XNOR2_X1 _15519_ (.A(_06393_),
    .B(\u0.subword[3] ),
    .ZN(_06394_));
 XNOR2_X1 _15520_ (.A(_06392_),
    .B(_06394_),
    .ZN(_06395_));
 MUX2_X1 _15521_ (.A(_06389_),
    .B(_06391_),
    .S(_06395_),
    .Z(_06396_));
 BUF_X8 _15522_ (.A(_06396_),
    .Z(_06397_));
 NAND2_X2 _15523_ (.A1(_06385_),
    .A2(_06397_),
    .ZN(_06398_));
 INV_X4 _15524_ (.A(_06398_),
    .ZN(_06399_));
 CLKBUF_X3 _15525_ (.A(_06399_),
    .Z(_06400_));
 BUF_X4 _15526_ (.A(_06400_),
    .Z(_00400_));
 BUF_X4 _15527_ (.A(_06279_),
    .Z(_06401_));
 AND2_X1 _15528_ (.A1(_06401_),
    .A2(net132),
    .ZN(_06402_));
 CLKBUF_X3 _15529_ (.A(\u0.w[0][4] ),
    .Z(_06403_));
 CLKBUF_X3 _15530_ (.A(\u0.w[1][4] ),
    .Z(_06404_));
 XNOR2_X2 _15531_ (.A(_06403_),
    .B(_06404_),
    .ZN(_06405_));
 CLKBUF_X3 _15532_ (.A(\u0.w[2][4] ),
    .Z(_06406_));
 CLKBUF_X3 _15533_ (.A(\u0.tmp_w[4] ),
    .Z(_06407_));
 XNOR2_X1 _15534_ (.A(_06407_),
    .B(\u0.subword[4] ),
    .ZN(_06408_));
 XNOR2_X1 _15535_ (.A(_06406_),
    .B(_06408_),
    .ZN(_06409_));
 XNOR2_X2 _15536_ (.A(_06405_),
    .B(_06409_),
    .ZN(_06410_));
 AOI21_X4 _15537_ (.A(_06402_),
    .B1(_06410_),
    .B2(_06267_),
    .ZN(_06411_));
 INV_X2 _15538_ (.A(_06411_),
    .ZN(_06412_));
 BUF_X4 _15539_ (.A(_06412_),
    .Z(_06413_));
 BUF_X4 _15540_ (.A(_06413_),
    .Z(_06414_));
 CLKBUF_X3 _15541_ (.A(_06414_),
    .Z(_00401_));
 INV_X1 _15542_ (.A(net163),
    .ZN(_06415_));
 CLKBUF_X3 _15543_ (.A(\u0.tmp_w[5] ),
    .Z(_06416_));
 CLKBUF_X3 _15544_ (.A(\u0.w[0][5] ),
    .Z(_06417_));
 CLKBUF_X3 _15545_ (.A(\u0.w[1][5] ),
    .Z(_06418_));
 XOR2_X2 _15546_ (.A(_06417_),
    .B(_06418_),
    .Z(_06419_));
 CLKBUF_X3 _15547_ (.A(\u0.w[2][5] ),
    .Z(_06420_));
 XNOR2_X1 _15548_ (.A(_06420_),
    .B(\u0.subword[5] ),
    .ZN(_06421_));
 XNOR2_X2 _15549_ (.A(_06419_),
    .B(_06421_),
    .ZN(_06422_));
 XNOR2_X1 _15550_ (.A(_06416_),
    .B(_06422_),
    .ZN(_06423_));
 MUX2_X1 _15551_ (.A(_06415_),
    .B(_06423_),
    .S(_06266_),
    .Z(_06424_));
 BUF_X4 _15552_ (.A(_06424_),
    .Z(_06425_));
 INV_X2 _15553_ (.A(_06425_),
    .ZN(_06426_));
 BUF_X4 _15554_ (.A(_06426_),
    .Z(_06427_));
 CLKBUF_X3 _15555_ (.A(_06427_),
    .Z(_00402_));
 BUF_X8 _15556_ (.A(_06267_),
    .Z(_06428_));
 NOR2_X1 _15557_ (.A1(_06428_),
    .A2(net183),
    .ZN(_06429_));
 BUF_X2 _15558_ (.A(\u0.tmp_w[6] ),
    .Z(_06430_));
 CLKBUF_X3 _15559_ (.A(\u0.w[0][6] ),
    .Z(_06431_));
 CLKBUF_X3 _15560_ (.A(\u0.w[1][6] ),
    .Z(_06432_));
 XOR2_X2 _15561_ (.A(_06431_),
    .B(_06432_),
    .Z(_06433_));
 BUF_X4 _15562_ (.A(\u0.w[2][6] ),
    .Z(_06434_));
 XNOR2_X1 _15563_ (.A(_06434_),
    .B(\u0.subword[6] ),
    .ZN(_06435_));
 XNOR2_X2 _15564_ (.A(_06433_),
    .B(_06435_),
    .ZN(_06436_));
 XNOR2_X2 _15565_ (.A(_06430_),
    .B(_06436_),
    .ZN(_06437_));
 AOI21_X4 _15566_ (.A(_06429_),
    .B1(_06437_),
    .B2(_06428_),
    .ZN(_06438_));
 BUF_X4 _15567_ (.A(_06438_),
    .Z(_00403_));
 CLKBUF_X3 _15568_ (.A(\u0.w[0][7] ),
    .Z(_06439_));
 CLKBUF_X3 _15569_ (.A(\u0.w[1][7] ),
    .Z(_06440_));
 XOR2_X2 _15570_ (.A(_06439_),
    .B(_06440_),
    .Z(_06441_));
 BUF_X4 _15571_ (.A(\u0.w[2][7] ),
    .Z(_06442_));
 XOR2_X2 _15572_ (.A(_06442_),
    .B(\u0.subword[7] ),
    .Z(_06443_));
 XNOR2_X2 _15573_ (.A(_06441_),
    .B(_06443_),
    .ZN(_06444_));
 XNOR2_X1 _15574_ (.A(\u0.tmp_w[7] ),
    .B(_06444_),
    .ZN(_06445_));
 MUX2_X1 _15575_ (.A(net201),
    .B(_06445_),
    .S(_06267_),
    .Z(_06446_));
 BUF_X4 _15576_ (.A(_06446_),
    .Z(_06447_));
 CLKBUF_X3 _15577_ (.A(_06447_),
    .Z(_06448_));
 CLKBUF_X3 _15578_ (.A(_06448_),
    .Z(_00404_));
 NOR2_X4 _15579_ (.A1(_06239_),
    .A2(net214),
    .ZN(_06449_));
 BUF_X4 _15580_ (.A(\u0.w[0][8] ),
    .Z(_06450_));
 BUF_X4 _15581_ (.A(\u0.w[1][8] ),
    .Z(_06451_));
 XOR2_X2 _15582_ (.A(_06450_),
    .B(_06451_),
    .Z(_06452_));
 NOR2_X1 _15583_ (.A1(_06339_),
    .A2(_06452_),
    .ZN(_06453_));
 XNOR2_X2 _15584_ (.A(_06450_),
    .B(_06451_),
    .ZN(_06454_));
 NOR2_X1 _15585_ (.A1(_06339_),
    .A2(_06454_),
    .ZN(_06455_));
 BUF_X4 _15586_ (.A(\u0.w[2][8] ),
    .Z(_06456_));
 BUF_X8 _15587_ (.A(\u0.tmp_w[8] ),
    .Z(_06457_));
 XNOR2_X2 _15588_ (.A(_06457_),
    .B(\u0.subword[8] ),
    .ZN(_06458_));
 XNOR2_X2 _15589_ (.A(_06456_),
    .B(_06458_),
    .ZN(_06459_));
 MUX2_X2 _15590_ (.A(_06453_),
    .B(_06455_),
    .S(_06459_),
    .Z(_06460_));
 NOR2_X4 _15591_ (.A1(_06449_),
    .A2(_06460_),
    .ZN(_06461_));
 INV_X2 _15592_ (.A(_06461_),
    .ZN(_06462_));
 BUF_X4 _15593_ (.A(_06462_),
    .Z(_06463_));
 BUF_X8 _15594_ (.A(_06463_),
    .Z(_14698_));
 NOR2_X1 _15595_ (.A1(_06239_),
    .A2(net225),
    .ZN(_06464_));
 BUF_X4 _15596_ (.A(\u0.w[0][9] ),
    .Z(_06465_));
 CLKBUF_X3 _15597_ (.A(\u0.w[1][9] ),
    .Z(_06466_));
 XNOR2_X2 _15598_ (.A(_06465_),
    .B(_06466_),
    .ZN(_06467_));
 AND2_X1 _15599_ (.A1(_06218_),
    .A2(_06467_),
    .ZN(_06468_));
 NOR2_X1 _15600_ (.A1(_06339_),
    .A2(_06467_),
    .ZN(_06469_));
 CLKBUF_X3 _15601_ (.A(\u0.w[2][9] ),
    .Z(_06470_));
 BUF_X1 rebuffer585 (.A(\u0.tmp_w[9] ),
    .Z(net1048));
 XNOR2_X2 _15603_ (.A(\u0.subword[9] ),
    .B(\u0.tmp_w[9] ),
    .ZN(_06472_));
 XNOR2_X2 _15604_ (.A(_06472_),
    .B(_06470_),
    .ZN(_06473_));
 MUX2_X2 _15605_ (.A(_06468_),
    .B(_06469_),
    .S(_06473_),
    .Z(_06474_));
 NOR2_X4 _15606_ (.A1(_06474_),
    .A2(_06464_),
    .ZN(_06475_));
 INV_X1 _15607_ (.A(net1233),
    .ZN(_06476_));
 BUF_X4 _15608_ (.A(_06476_),
    .Z(_06477_));
 BUF_X8 _15609_ (.A(_06477_),
    .Z(_14703_));
 NAND2_X1 _15610_ (.A1(_06245_),
    .A2(net34),
    .ZN(_06478_));
 CLKBUF_X3 _15611_ (.A(\u0.tmp_w[10] ),
    .Z(_06479_));
 BUF_X4 _15612_ (.A(\u0.w[0][10] ),
    .Z(_06480_));
 XOR2_X2 _15613_ (.A(_06480_),
    .B(_00410_),
    .Z(_06481_));
 BUF_X4 _15614_ (.A(\u0.w[2][10] ),
    .Z(_06482_));
 BUF_X4 _15615_ (.A(\u0.w[1][10] ),
    .Z(_06483_));
 NOR2_X1 _15616_ (.A1(_06482_),
    .A2(_06483_),
    .ZN(_06484_));
 NAND4_X1 _15617_ (.A1(_06220_),
    .A2(_06479_),
    .A3(_06481_),
    .A4(_06484_),
    .ZN(_06485_));
 INV_X1 _15618_ (.A(_06483_),
    .ZN(_06486_));
 NOR2_X1 _15619_ (.A1(_06216_),
    .A2(_06479_),
    .ZN(_06487_));
 NAND4_X1 _15620_ (.A1(_06482_),
    .A2(_06486_),
    .A3(_06481_),
    .A4(_06487_),
    .ZN(_06488_));
 INV_X1 _15621_ (.A(_06482_),
    .ZN(_06489_));
 NAND4_X1 _15622_ (.A1(_06489_),
    .A2(_06483_),
    .A3(_06481_),
    .A4(_06487_),
    .ZN(_06490_));
 INV_X2 _15623_ (.A(_06479_),
    .ZN(_06491_));
 XNOR2_X2 _15624_ (.A(_06480_),
    .B(_00410_),
    .ZN(_06492_));
 NAND2_X1 _15625_ (.A1(\u0.w[2][10] ),
    .A2(\u0.w[1][10] ),
    .ZN(_06493_));
 OR4_X1 _15626_ (.A1(_06216_),
    .A2(_06491_),
    .A3(_06492_),
    .A4(_06493_),
    .ZN(_06494_));
 AND4_X1 _15627_ (.A1(_06485_),
    .A2(_06488_),
    .A3(_06490_),
    .A4(_06494_),
    .ZN(_06495_));
 AND2_X1 _15628_ (.A1(_06484_),
    .A2(_06487_),
    .ZN(_06496_));
 NOR4_X1 _15629_ (.A1(_06226_),
    .A2(_06491_),
    .A3(_06489_),
    .A4(_06483_),
    .ZN(_06497_));
 OAI21_X1 _15630_ (.A(_06492_),
    .B1(_06496_),
    .B2(_06497_),
    .ZN(_06498_));
 NOR4_X1 _15631_ (.A1(_06226_),
    .A2(_06491_),
    .A3(_06482_),
    .A4(_06486_),
    .ZN(_06499_));
 NOR3_X1 _15632_ (.A1(net16),
    .A2(_06479_),
    .A3(_06493_),
    .ZN(_06500_));
 OAI21_X1 _15633_ (.A(_06492_),
    .B1(_06499_),
    .B2(_06500_),
    .ZN(_06501_));
 AND4_X4 _15634_ (.A1(_06478_),
    .A2(_06495_),
    .A3(_06498_),
    .A4(_06501_),
    .ZN(_06502_));
 BUF_X8 _15635_ (.A(_06502_),
    .Z(_06503_));
 INV_X4 _15636_ (.A(_06503_),
    .ZN(_06504_));
 BUF_X8 _15637_ (.A(_06504_),
    .Z(_06505_));
 BUF_X4 _15638_ (.A(_06505_),
    .Z(_06506_));
 BUF_X4 _15639_ (.A(_06506_),
    .Z(_06507_));
 BUF_X8 _15640_ (.A(_06507_),
    .Z(_14717_));
 OR2_X1 _15641_ (.A1(_06218_),
    .A2(net52),
    .ZN(_06508_));
 BUF_X8 _15642_ (.A(_06508_),
    .Z(_06509_));
 BUF_X4 _15643_ (.A(\u0.w[0][11] ),
    .Z(_06510_));
 BUF_X4 _15644_ (.A(\u0.w[1][11] ),
    .Z(_06511_));
 XNOR2_X2 _15645_ (.A(_06510_),
    .B(_06511_),
    .ZN(_06512_));
 NAND2_X1 _15646_ (.A1(_06217_),
    .A2(_06512_),
    .ZN(_06513_));
 XOR2_X2 _15647_ (.A(_06510_),
    .B(_06511_),
    .Z(_06514_));
 NAND2_X1 _15648_ (.A1(_06217_),
    .A2(_06514_),
    .ZN(_06515_));
 BUF_X4 _15649_ (.A(\u0.w[2][11] ),
    .Z(_06516_));
 BUF_X4 _15650_ (.A(\u0.tmp_w[11] ),
    .Z(_06517_));
 XNOR2_X1 _15651_ (.A(_06517_),
    .B(\u0.subword[11] ),
    .ZN(_06518_));
 XNOR2_X1 _15652_ (.A(_06516_),
    .B(_06518_),
    .ZN(_06519_));
 MUX2_X2 _15653_ (.A(_06513_),
    .B(_06515_),
    .S(_06519_),
    .Z(_06520_));
 BUF_X8 _15654_ (.A(_06520_),
    .Z(_06521_));
 NAND2_X4 _15655_ (.A1(_06509_),
    .A2(_06521_),
    .ZN(_06522_));
 INV_X2 _15656_ (.A(_06522_),
    .ZN(_06523_));
 BUF_X4 _15657_ (.A(_06523_),
    .Z(_06524_));
 CLKBUF_X3 _15658_ (.A(_06524_),
    .Z(_06525_));
 BUF_X4 _15659_ (.A(_06525_),
    .Z(_00385_));
 NOR2_X1 _15660_ (.A1(_06239_),
    .A2(net62),
    .ZN(_06526_));
 CLKBUF_X3 _15661_ (.A(\u0.w[0][12] ),
    .Z(_06527_));
 CLKBUF_X3 _15662_ (.A(\u0.w[1][12] ),
    .Z(_06528_));
 XNOR2_X2 _15663_ (.A(_06527_),
    .B(_06528_),
    .ZN(_06529_));
 AND2_X1 _15664_ (.A1(_06218_),
    .A2(_06529_),
    .ZN(_06530_));
 NOR2_X1 _15665_ (.A1(_06245_),
    .A2(_06529_),
    .ZN(_06531_));
 BUF_X4 _15666_ (.A(\u0.w[2][12] ),
    .Z(_06532_));
 CLKBUF_X3 _15667_ (.A(\u0.tmp_w[12] ),
    .Z(_06533_));
 XNOR2_X1 _15668_ (.A(_06533_),
    .B(\u0.subword[12] ),
    .ZN(_06534_));
 XNOR2_X1 _15669_ (.A(_06532_),
    .B(_06534_),
    .ZN(_06535_));
 MUX2_X1 _15670_ (.A(_06530_),
    .B(_06531_),
    .S(_06535_),
    .Z(_06536_));
 OR2_X1 _15671_ (.A1(_06526_),
    .A2(_06536_),
    .ZN(_06537_));
 INV_X2 _15672_ (.A(_06537_),
    .ZN(_06538_));
 BUF_X4 _15673_ (.A(_06538_),
    .Z(_06539_));
 BUF_X4 _15674_ (.A(_06539_),
    .Z(_06540_));
 BUF_X4 _15675_ (.A(_06540_),
    .Z(_00386_));
 INV_X1 _15676_ (.A(net63),
    .ZN(_06541_));
 CLKBUF_X3 _15677_ (.A(\u0.w[0][13] ),
    .Z(_06542_));
 CLKBUF_X3 _15678_ (.A(\u0.w[1][13] ),
    .Z(_06543_));
 XNOR2_X1 _15679_ (.A(_06542_),
    .B(_06543_),
    .ZN(_06544_));
 BUF_X4 _15680_ (.A(\u0.w[2][13] ),
    .Z(_06545_));
 BUF_X4 _15681_ (.A(\u0.tmp_w[13] ),
    .Z(_06546_));
 XOR2_X1 _15682_ (.A(_06546_),
    .B(\u0.subword[13] ),
    .Z(_06547_));
 XNOR2_X1 _15683_ (.A(_06545_),
    .B(_06547_),
    .ZN(_06548_));
 XNOR2_X1 _15684_ (.A(_06544_),
    .B(_06548_),
    .ZN(_06549_));
 MUX2_X2 _15685_ (.A(_06541_),
    .B(_06549_),
    .S(_06266_),
    .Z(_06550_));
 INV_X4 _15686_ (.A(_06550_),
    .ZN(_06551_));
 CLKBUF_X3 _15687_ (.A(_06551_),
    .Z(_06552_));
 CLKBUF_X3 _15688_ (.A(_06552_),
    .Z(_00387_));
 NOR2_X1 _15689_ (.A1(_06428_),
    .A2(net67),
    .ZN(_06553_));
 CLKBUF_X3 _15690_ (.A(\u0.tmp_w[14] ),
    .Z(_06554_));
 BUF_X4 _15691_ (.A(\u0.w[0][14] ),
    .Z(_06555_));
 BUF_X2 _15692_ (.A(\u0.w[1][14] ),
    .Z(_06556_));
 XOR2_X2 _15693_ (.A(_06555_),
    .B(_06556_),
    .Z(_06557_));
 BUF_X4 _15694_ (.A(\u0.w[2][14] ),
    .Z(_06558_));
 XNOR2_X1 _15695_ (.A(_06558_),
    .B(\u0.subword[14] ),
    .ZN(_06559_));
 XNOR2_X2 _15696_ (.A(_06557_),
    .B(_06559_),
    .ZN(_06560_));
 XNOR2_X2 _15697_ (.A(_06554_),
    .B(_06560_),
    .ZN(_06561_));
 AOI21_X4 _15698_ (.A(_06553_),
    .B1(_06561_),
    .B2(_06428_),
    .ZN(_06562_));
 BUF_X4 _15699_ (.A(_06562_),
    .Z(_00388_));
 CLKBUF_X3 _15700_ (.A(\u0.tmp_w[15] ),
    .Z(_06563_));
 BUF_X2 _15701_ (.A(\u0.w[0][15] ),
    .Z(_06564_));
 CLKBUF_X3 _15702_ (.A(\u0.w[1][15] ),
    .Z(_06565_));
 XOR2_X2 _15703_ (.A(_06564_),
    .B(_06565_),
    .Z(_06566_));
 BUF_X4 _15704_ (.A(\u0.w[2][15] ),
    .Z(_06567_));
 XNOR2_X1 _15705_ (.A(_06567_),
    .B(\u0.subword[15] ),
    .ZN(_06568_));
 XNOR2_X2 _15706_ (.A(_06566_),
    .B(_06568_),
    .ZN(_06569_));
 XNOR2_X1 _15707_ (.A(_06563_),
    .B(_06569_),
    .ZN(_06570_));
 NAND2_X1 _15708_ (.A1(_06266_),
    .A2(_06570_),
    .ZN(_06571_));
 OAI21_X4 _15709_ (.A(_06571_),
    .B1(net68),
    .B2(_06267_),
    .ZN(_06572_));
 INV_X4 _15710_ (.A(_06572_),
    .ZN(_06573_));
 CLKBUF_X3 _15711_ (.A(_06573_),
    .Z(_00389_));
 CLKBUF_X3 _15712_ (.A(\u0.tmp_w[22] ),
    .Z(_06574_));
 CLKBUF_X3 _15713_ (.A(\u0.w[0][22] ),
    .Z(_06575_));
 BUF_X4 _15714_ (.A(\u0.w[1][22] ),
    .Z(_06576_));
 XOR2_X2 _15715_ (.A(_06575_),
    .B(_06576_),
    .Z(_06577_));
 BUF_X4 _15716_ (.A(\u0.w[2][22] ),
    .Z(_06578_));
 XNOR2_X1 _15717_ (.A(_06578_),
    .B(\u0.subword[22] ),
    .ZN(_06579_));
 XNOR2_X1 _15718_ (.A(_06577_),
    .B(_06579_),
    .ZN(_06580_));
 XNOR2_X1 _15719_ (.A(_06574_),
    .B(_06580_),
    .ZN(_06581_));
 NAND2_X1 _15720_ (.A1(_06428_),
    .A2(_06581_),
    .ZN(_06582_));
 OAI21_X4 _15721_ (.A(_06582_),
    .B1(net77),
    .B2(_06428_),
    .ZN(_06583_));
 INV_X1 _15722_ (.A(_06583_),
    .ZN(_06584_));
 BUF_X4 _15723_ (.A(_06584_),
    .Z(_06585_));
 CLKBUF_X3 _15724_ (.A(_06585_),
    .Z(_00393_));
 CLKBUF_X3 _15725_ (.A(\u0.tmp_w[23] ),
    .Z(_06586_));
 BUF_X4 _15726_ (.A(\u0.w[0][23] ),
    .Z(_06587_));
 BUF_X4 _15727_ (.A(\u0.w[1][23] ),
    .Z(_06588_));
 XOR2_X2 _15728_ (.A(_06587_),
    .B(_06588_),
    .Z(_06589_));
 BUF_X4 _15729_ (.A(\u0.w[2][23] ),
    .Z(_06590_));
 XNOR2_X1 _15730_ (.A(_06590_),
    .B(\u0.subword[23] ),
    .ZN(_06591_));
 XNOR2_X1 _15731_ (.A(_06589_),
    .B(_06591_),
    .ZN(_06592_));
 XNOR2_X1 _15732_ (.A(_06586_),
    .B(_06592_),
    .ZN(_06593_));
 NAND2_X1 _15733_ (.A1(_06267_),
    .A2(_06593_),
    .ZN(_06594_));
 OAI21_X2 _15734_ (.A(_06594_),
    .B1(net78),
    .B2(_06267_),
    .ZN(_06595_));
 INV_X2 _15735_ (.A(_06595_),
    .ZN(_06596_));
 BUF_X4 _15736_ (.A(_06596_),
    .Z(_00394_));
 AND2_X2 _15737_ (.A1(_06279_),
    .A2(net79),
    .ZN(_06597_));
 CLKBUF_X3 _15738_ (.A(\u0.w[0][24] ),
    .Z(_06598_));
 XNOR2_X2 _15739_ (.A(_06598_),
    .B(\u0.subword[24] ),
    .ZN(_06599_));
 AND2_X1 _15740_ (.A1(_06220_),
    .A2(_06599_),
    .ZN(_06600_));
 NOR2_X1 _15741_ (.A1(_06245_),
    .A2(_06599_),
    .ZN(_06601_));
 BUF_X1 rebuffer323 (.A(\u0.tmp_w[24] ),
    .Z(net786));
 XNOR2_X2 _15743_ (.A(\u0.tmp_w[24] ),
    .B(\u0.r0.out[24] ),
    .ZN(_06603_));
 BUF_X4 _15744_ (.A(\u0.w[2][24] ),
    .Z(_06604_));
 BUF_X1 rebuffer319 (.A(\u0.w[1][24] ),
    .Z(net782));
 XNOR2_X2 _15746_ (.A(_06604_),
    .B(\u0.w[1][24] ),
    .ZN(_06606_));
 XNOR2_X2 _15747_ (.A(_06603_),
    .B(_06606_),
    .ZN(_06607_));
 MUX2_X2 _15748_ (.A(_06600_),
    .B(_06601_),
    .S(_06607_),
    .Z(_06608_));
 OR2_X4 _15749_ (.A1(_06608_),
    .A2(_06597_),
    .ZN(_06609_));
 BUF_X16 _15750_ (.A(_06609_),
    .Z(_06610_));
 INV_X32 _15751_ (.A(_06610_),
    .ZN(_06611_));
 BUF_X32 _15752_ (.A(_06611_),
    .Z(_06612_));
 BUF_X32 _15753_ (.A(_06612_),
    .Z(_14766_));
 NAND2_X2 _15754_ (.A1(_06279_),
    .A2(net80),
    .ZN(_06613_));
 BUF_X4 _15755_ (.A(\u0.w[0][25] ),
    .Z(_06614_));
 XNOR2_X2 _15756_ (.A(_06614_),
    .B(\u0.subword[25] ),
    .ZN(_06615_));
 NAND2_X1 _15757_ (.A1(_06218_),
    .A2(_06615_),
    .ZN(_06616_));
 XOR2_X2 _15758_ (.A(_06614_),
    .B(\u0.subword[25] ),
    .Z(_06617_));
 NAND2_X1 _15759_ (.A1(_06218_),
    .A2(_06617_),
    .ZN(_06618_));
 BUF_X4 _15760_ (.A(\u0.tmp_w[25] ),
    .Z(_06619_));
 XNOR2_X1 _15761_ (.A(_06619_),
    .B(\u0.r0.out[25] ),
    .ZN(_06620_));
 BUF_X1 rebuffer332 (.A(\u0.tmp_w[24] ),
    .Z(net795));
 BUF_X1 rebuffer624 (.A(\u0.w[1][25] ),
    .Z(net1087));
 XNOR2_X2 _15764_ (.A(\u0.w[1][25] ),
    .B(\u0.w[2][25] ),
    .ZN(_06623_));
 XNOR2_X2 _15765_ (.A(_06620_),
    .B(_06623_),
    .ZN(_06624_));
 MUX2_X2 _15766_ (.A(_06616_),
    .B(_06618_),
    .S(_06624_),
    .Z(_06625_));
 NAND2_X4 _15767_ (.A1(_06613_),
    .A2(_06625_),
    .ZN(_06626_));
 INV_X2 _15768_ (.A(_06626_),
    .ZN(_06627_));
 BUF_X8 _15769_ (.A(_06627_),
    .Z(_06628_));
 BUF_X8 _15770_ (.A(_06628_),
    .Z(_14771_));
 NAND2_X2 _15771_ (.A1(net18),
    .A2(net81),
    .ZN(_06629_));
 BUF_X4 _15772_ (.A(\u0.w[0][26] ),
    .Z(_06630_));
 XNOR2_X2 _15773_ (.A(_06630_),
    .B(\u0.subword[26] ),
    .ZN(_06631_));
 NAND2_X1 _15774_ (.A1(_06220_),
    .A2(_06631_),
    .ZN(_06632_));
 XOR2_X2 _15775_ (.A(_06630_),
    .B(\u0.subword[26] ),
    .Z(_06633_));
 NAND2_X1 _15776_ (.A1(_06220_),
    .A2(_06633_),
    .ZN(_06634_));
 BUF_X2 _15777_ (.A(\u0.tmp_w[26] ),
    .Z(_06635_));
 XNOR2_X1 _15778_ (.A(_06635_),
    .B(\u0.r0.out[26] ),
    .ZN(_06636_));
 CLKBUF_X3 _15779_ (.A(\u0.w[2][26] ),
    .Z(_06637_));
 BUF_X4 _15780_ (.A(\u0.w[1][26] ),
    .Z(_06638_));
 XNOR2_X2 _15781_ (.A(_06637_),
    .B(_06638_),
    .ZN(_06639_));
 XNOR2_X2 _15782_ (.A(_06636_),
    .B(_06639_),
    .ZN(_06640_));
 MUX2_X2 _15783_ (.A(_06632_),
    .B(_06634_),
    .S(_06640_),
    .Z(_06641_));
 NAND2_X1 _15784_ (.A1(_06629_),
    .A2(_06641_),
    .ZN(_06642_));
 INV_X2 _15785_ (.A(_06642_),
    .ZN(_06643_));
 BUF_X4 _15786_ (.A(_06643_),
    .Z(_06644_));
 BUF_X4 _15787_ (.A(_06644_),
    .Z(_06645_));
 BUF_X4 _15788_ (.A(_06645_),
    .Z(_14785_));
 BUF_X2 _15789_ (.A(key[27]),
    .Z(_06646_));
 AND2_X4 _15790_ (.A1(net18),
    .A2(_06646_),
    .ZN(_06647_));
 BUF_X8 _15791_ (.A(_06647_),
    .Z(_06648_));
 BUF_X4 _15792_ (.A(\u0.w[0][27] ),
    .Z(_06649_));
 XOR2_X2 _15793_ (.A(_06649_),
    .B(\u0.subword[27] ),
    .Z(_06650_));
 NOR2_X1 _15794_ (.A1(net6),
    .A2(_06650_),
    .ZN(_06651_));
 XNOR2_X2 _15795_ (.A(_06649_),
    .B(\u0.subword[27] ),
    .ZN(_06652_));
 NOR2_X1 _15796_ (.A1(net6),
    .A2(_06652_),
    .ZN(_06653_));
 BUF_X2 _15797_ (.A(\u0.tmp_w[27] ),
    .Z(_06654_));
 XNOR2_X1 _15798_ (.A(_06654_),
    .B(\u0.r0.out[27] ),
    .ZN(_06655_));
 BUF_X2 _15799_ (.A(\u0.w[2][27] ),
    .Z(_06656_));
 CLKBUF_X3 _15800_ (.A(\u0.w[1][27] ),
    .Z(_06657_));
 XNOR2_X2 _15801_ (.A(_06656_),
    .B(_06657_),
    .ZN(_06658_));
 XNOR2_X1 _15802_ (.A(_06655_),
    .B(_06658_),
    .ZN(_06659_));
 MUX2_X1 _15803_ (.A(_06651_),
    .B(_06653_),
    .S(_06659_),
    .Z(_06660_));
 BUF_X4 _15804_ (.A(_06660_),
    .Z(_06661_));
 NOR2_X4 _15805_ (.A1(_06648_),
    .A2(_06661_),
    .ZN(_06662_));
 INV_X4 _15806_ (.A(_06662_),
    .ZN(_06663_));
 BUF_X4 _15807_ (.A(_06663_),
    .Z(_06664_));
 BUF_X4 _15808_ (.A(_06664_),
    .Z(_00395_));
 AND2_X1 _15809_ (.A1(_06401_),
    .A2(net82),
    .ZN(_06665_));
 CLKBUF_X3 _15810_ (.A(\u0.w[0][28] ),
    .Z(_06666_));
 XNOR2_X2 _15811_ (.A(_06666_),
    .B(\u0.subword[28] ),
    .ZN(_06667_));
 AND2_X1 _15812_ (.A1(_06239_),
    .A2(_06667_),
    .ZN(_06668_));
 NOR2_X1 _15813_ (.A1(_06279_),
    .A2(_06667_),
    .ZN(_06669_));
 CLKBUF_X3 _15814_ (.A(\u0.tmp_w[28] ),
    .Z(_06670_));
 XNOR2_X1 _15815_ (.A(_06670_),
    .B(\u0.r0.out[28] ),
    .ZN(_06671_));
 CLKBUF_X3 _15816_ (.A(\u0.w[2][28] ),
    .Z(_06672_));
 BUF_X2 _15817_ (.A(\u0.w[1][28] ),
    .Z(_06673_));
 XNOR2_X2 _15818_ (.A(_06672_),
    .B(_06673_),
    .ZN(_06674_));
 XNOR2_X1 _15819_ (.A(_06671_),
    .B(_06674_),
    .ZN(_06675_));
 MUX2_X2 _15820_ (.A(_06668_),
    .B(_06669_),
    .S(_06675_),
    .Z(_06676_));
 NOR2_X4 _15821_ (.A1(_06665_),
    .A2(_06676_),
    .ZN(_06677_));
 INV_X2 _15822_ (.A(_06677_),
    .ZN(_06678_));
 BUF_X4 _15823_ (.A(_06678_),
    .Z(_06679_));
 BUF_X4 _15824_ (.A(_06679_),
    .Z(_06680_));
 BUF_X4 _15825_ (.A(_06680_),
    .Z(_06681_));
 CLKBUF_X3 _15826_ (.A(_06681_),
    .Z(_00396_));
 AND2_X1 _15827_ (.A1(_06279_),
    .A2(net83),
    .ZN(_06682_));
 CLKBUF_X3 _15828_ (.A(\u0.w[0][29] ),
    .Z(_06683_));
 XOR2_X2 _15829_ (.A(_06683_),
    .B(\u0.subword[29] ),
    .Z(_06684_));
 CLKBUF_X3 _15830_ (.A(\u0.tmp_w[29] ),
    .Z(_06685_));
 XNOR2_X1 _15831_ (.A(_06685_),
    .B(\u0.r0.out[29] ),
    .ZN(_06686_));
 CLKBUF_X3 _15832_ (.A(\u0.w[2][29] ),
    .Z(_06687_));
 CLKBUF_X3 _15833_ (.A(\u0.w[1][29] ),
    .Z(_06688_));
 XNOR2_X2 _15834_ (.A(_06687_),
    .B(_06688_),
    .ZN(_06689_));
 XNOR2_X1 _15835_ (.A(_06686_),
    .B(_06689_),
    .ZN(_06690_));
 XNOR2_X2 _15836_ (.A(_06684_),
    .B(_06690_),
    .ZN(_06691_));
 AOI21_X4 _15837_ (.A(_06682_),
    .B1(_06691_),
    .B2(_06266_),
    .ZN(_06692_));
 INV_X1 _15838_ (.A(_06692_),
    .ZN(_06693_));
 BUF_X4 _15839_ (.A(_06693_),
    .Z(_06694_));
 CLKBUF_X3 _15840_ (.A(_06694_),
    .Z(_06695_));
 CLKBUF_X3 _15841_ (.A(_06695_),
    .Z(_00397_));
 BUF_X2 _15842_ (.A(\u0.w[2][30] ),
    .Z(_06696_));
 CLKBUF_X3 _15843_ (.A(\u0.w[1][30] ),
    .Z(_06697_));
 XOR2_X2 _15844_ (.A(_06696_),
    .B(_06697_),
    .Z(_06698_));
 BUF_X2 _15845_ (.A(\u0.tmp_w[30] ),
    .Z(_06699_));
 XNOR2_X1 _15846_ (.A(_06699_),
    .B(\u0.r0.out[30] ),
    .ZN(_06700_));
 CLKBUF_X3 _15847_ (.A(\u0.w[0][30] ),
    .Z(_06701_));
 XNOR2_X2 _15848_ (.A(_06701_),
    .B(\u0.subword[30] ),
    .ZN(_06702_));
 XNOR2_X1 _15849_ (.A(_06700_),
    .B(_06702_),
    .ZN(_06703_));
 XNOR2_X1 _15850_ (.A(_06698_),
    .B(_06703_),
    .ZN(_06704_));
 MUX2_X1 _15851_ (.A(net85),
    .B(_06704_),
    .S(_06428_),
    .Z(_06705_));
 BUF_X4 _15852_ (.A(_06705_),
    .Z(_00398_));
 CLKBUF_X3 _15853_ (.A(\u0.w[0][31] ),
    .Z(_06706_));
 XNOR2_X2 _15854_ (.A(_06706_),
    .B(\u0.subword[31] ),
    .ZN(_06707_));
 CLKBUF_X3 _15855_ (.A(\u0.tmp_w[31] ),
    .Z(_06708_));
 XNOR2_X1 _15856_ (.A(_06708_),
    .B(\u0.r0.out[31] ),
    .ZN(_06709_));
 CLKBUF_X3 _15857_ (.A(\u0.w[2][31] ),
    .Z(_06710_));
 BUF_X2 _15858_ (.A(\u0.w[1][31] ),
    .Z(_06711_));
 XNOR2_X2 _15859_ (.A(_06710_),
    .B(_06711_),
    .ZN(_06712_));
 XNOR2_X1 _15860_ (.A(_06709_),
    .B(_06712_),
    .ZN(_06713_));
 XNOR2_X1 _15861_ (.A(_06707_),
    .B(_06713_),
    .ZN(_06714_));
 NAND2_X1 _15862_ (.A1(_06428_),
    .A2(_06714_),
    .ZN(_06715_));
 OAI21_X4 _15863_ (.A(_06715_),
    .B1(net86),
    .B2(_06428_),
    .ZN(_06716_));
 INV_X1 _15864_ (.A(_06716_),
    .ZN(_06717_));
 BUF_X4 _15865_ (.A(_06717_),
    .Z(_00399_));
 XNOR2_X1 _15866_ (.A(_00411_),
    .B(_06327_),
    .ZN(_06718_));
 XNOR2_X1 _15867_ (.A(_06330_),
    .B(_06718_),
    .ZN(_06719_));
 BUF_X4 _15868_ (.A(_06428_),
    .Z(_06720_));
 BUF_X4 _15869_ (.A(_06720_),
    .Z(_06721_));
 MUX2_X1 _15870_ (.A(net87),
    .B(_06719_),
    .S(_06721_),
    .Z(_00353_));
 XNOR2_X1 _15871_ (.A(_00412_),
    .B(_06344_),
    .ZN(_06722_));
 XNOR2_X1 _15872_ (.A(_06346_),
    .B(_06722_),
    .ZN(_06723_));
 MUX2_X1 _15873_ (.A(net88),
    .B(_06723_),
    .S(_06721_),
    .Z(_00364_));
 XNOR2_X1 _15874_ (.A(_06359_),
    .B(net1162),
    .ZN(_06724_));
 XNOR2_X1 _15875_ (.A(_06358_),
    .B(_06724_),
    .ZN(_06725_));
 BUF_X4 _15876_ (.A(_06720_),
    .Z(_06726_));
 MUX2_X1 _15877_ (.A(net89),
    .B(_06725_),
    .S(_06726_),
    .Z(_00375_));
 XNOR2_X1 _15878_ (.A(_00413_),
    .B(_06388_),
    .ZN(_06727_));
 XNOR2_X1 _15879_ (.A(_06392_),
    .B(_06727_),
    .ZN(_06728_));
 MUX2_X1 _15880_ (.A(net90),
    .B(_06728_),
    .S(_06726_),
    .Z(_00378_));
 XNOR2_X1 _15881_ (.A(_00414_),
    .B(_06405_),
    .ZN(_06729_));
 XNOR2_X1 _15882_ (.A(_06406_),
    .B(_06729_),
    .ZN(_06730_));
 MUX2_X1 _15883_ (.A(net91),
    .B(_06730_),
    .S(_06726_),
    .Z(_00379_));
 XOR2_X2 _15884_ (.A(_00415_),
    .B(_06419_),
    .Z(_06731_));
 XNOR2_X1 _15885_ (.A(_06420_),
    .B(_06731_),
    .ZN(_06732_));
 MUX2_X1 _15886_ (.A(net92),
    .B(_06732_),
    .S(_06726_),
    .Z(_00380_));
 XOR2_X2 _15887_ (.A(_00416_),
    .B(_06433_),
    .Z(_06733_));
 XNOR2_X1 _15888_ (.A(_06434_),
    .B(_06733_),
    .ZN(_06734_));
 MUX2_X1 _15889_ (.A(net104),
    .B(_06734_),
    .S(_06726_),
    .Z(_00381_));
 XOR2_X2 _15890_ (.A(_00417_),
    .B(_06441_),
    .Z(_06735_));
 XNOR2_X1 _15891_ (.A(_06442_),
    .B(_06735_),
    .ZN(_06736_));
 MUX2_X1 _15892_ (.A(net115),
    .B(_06736_),
    .S(_06726_),
    .Z(_00382_));
 XNOR2_X1 _15893_ (.A(_00418_),
    .B(_06454_),
    .ZN(_06737_));
 XNOR2_X1 _15894_ (.A(_06456_),
    .B(_06737_),
    .ZN(_06738_));
 MUX2_X1 _15895_ (.A(net117),
    .B(_06738_),
    .S(_06726_),
    .Z(_00383_));
 XNOR2_X1 _15896_ (.A(_00419_),
    .B(_06467_),
    .ZN(_06739_));
 XNOR2_X1 _15897_ (.A(_06470_),
    .B(_06739_),
    .ZN(_06740_));
 MUX2_X1 _15898_ (.A(net118),
    .B(_06740_),
    .S(_06726_),
    .Z(_00384_));
 XNOR2_X1 _15899_ (.A(_06483_),
    .B(_06492_),
    .ZN(_06741_));
 XNOR2_X1 _15900_ (.A(_06482_),
    .B(_06741_),
    .ZN(_06742_));
 MUX2_X1 _15901_ (.A(net119),
    .B(_06742_),
    .S(_06726_),
    .Z(_00354_));
 XNOR2_X1 _15902_ (.A(_00420_),
    .B(_06512_),
    .ZN(_06743_));
 XNOR2_X1 _15903_ (.A(_06516_),
    .B(_06743_),
    .ZN(_06744_));
 MUX2_X1 _15904_ (.A(net120),
    .B(_06744_),
    .S(_06726_),
    .Z(_00355_));
 XNOR2_X1 _15905_ (.A(_00421_),
    .B(_06529_),
    .ZN(_06745_));
 XNOR2_X1 _15906_ (.A(_06532_),
    .B(_06745_),
    .ZN(_06746_));
 BUF_X4 _15907_ (.A(_06720_),
    .Z(_06747_));
 MUX2_X1 _15908_ (.A(net121),
    .B(_06746_),
    .S(_06747_),
    .Z(_00356_));
 XNOR2_X1 _15909_ (.A(_00422_),
    .B(_06544_),
    .ZN(_06748_));
 XNOR2_X1 _15910_ (.A(_06545_),
    .B(_06748_),
    .ZN(_06749_));
 MUX2_X1 _15911_ (.A(net127),
    .B(_06749_),
    .S(_06747_),
    .Z(_00357_));
 XOR2_X2 _15912_ (.A(_00423_),
    .B(_06557_),
    .Z(_06750_));
 XNOR2_X1 _15913_ (.A(_06558_),
    .B(_06750_),
    .ZN(_06751_));
 MUX2_X1 _15914_ (.A(net128),
    .B(_06751_),
    .S(_06747_),
    .Z(_00358_));
 XOR2_X2 _15915_ (.A(_00424_),
    .B(_06566_),
    .Z(_06752_));
 XNOR2_X1 _15916_ (.A(_06567_),
    .B(_06752_),
    .ZN(_06753_));
 MUX2_X1 _15917_ (.A(net129),
    .B(_06753_),
    .S(_06747_),
    .Z(_00359_));
 XNOR2_X1 _15918_ (.A(_00425_),
    .B(_06243_),
    .ZN(_06754_));
 XNOR2_X1 _15919_ (.A(_06247_),
    .B(_06754_),
    .ZN(_06755_));
 MUX2_X1 _15920_ (.A(net130),
    .B(_06755_),
    .S(_06747_),
    .Z(_00360_));
 XNOR2_X1 _15921_ (.A(_00426_),
    .B(_06257_),
    .ZN(_06756_));
 XNOR2_X1 _15922_ (.A(_06260_),
    .B(_06756_),
    .ZN(_06757_));
 MUX2_X1 _15923_ (.A(net131),
    .B(_06757_),
    .S(_06747_),
    .Z(_00361_));
 XNOR2_X1 _15924_ (.A(_06303_),
    .B(_06309_),
    .ZN(_06758_));
 XNOR2_X1 _15925_ (.A(_06306_),
    .B(_06758_),
    .ZN(_06759_));
 MUX2_X1 _15926_ (.A(net134),
    .B(_06759_),
    .S(_06747_),
    .Z(_00362_));
 XNOR2_X1 _15927_ (.A(_00427_),
    .B(_06223_),
    .ZN(_06760_));
 XNOR2_X1 _15928_ (.A(_06228_),
    .B(_06760_),
    .ZN(_06761_));
 MUX2_X1 _15929_ (.A(net135),
    .B(_06761_),
    .S(_06747_),
    .Z(_00363_));
 XNOR2_X1 _15930_ (.A(_00428_),
    .B(_06283_),
    .ZN(_06762_));
 XNOR2_X1 _15931_ (.A(_06284_),
    .B(_06762_),
    .ZN(_06763_));
 MUX2_X1 _15932_ (.A(net136),
    .B(_06763_),
    .S(_06747_),
    .Z(_00365_));
 XOR2_X2 _15933_ (.A(_00429_),
    .B(_06271_),
    .Z(_06764_));
 XNOR2_X1 _15934_ (.A(_06272_),
    .B(_06764_),
    .ZN(_06765_));
 MUX2_X1 _15935_ (.A(net137),
    .B(_06765_),
    .S(_06747_),
    .Z(_00366_));
 XOR2_X2 _15936_ (.A(_00430_),
    .B(_06577_),
    .Z(_06766_));
 XNOR2_X1 _15937_ (.A(_06578_),
    .B(_06766_),
    .ZN(_06767_));
 BUF_X4 _15938_ (.A(_06720_),
    .Z(_06768_));
 MUX2_X1 _15939_ (.A(net142),
    .B(_06767_),
    .S(_06768_),
    .Z(_00367_));
 XOR2_X2 _15940_ (.A(_00431_),
    .B(_06589_),
    .Z(_06769_));
 XNOR2_X1 _15941_ (.A(_06590_),
    .B(_06769_),
    .ZN(_06770_));
 MUX2_X1 _15942_ (.A(net147),
    .B(_06770_),
    .S(_06768_),
    .Z(_00368_));
 BUF_X4 _15943_ (.A(_06401_),
    .Z(_06771_));
 BUF_X4 _15944_ (.A(_06771_),
    .Z(_06772_));
 NAND2_X1 _15945_ (.A1(_06772_),
    .A2(net148),
    .ZN(_06773_));
 XNOR2_X2 _15946_ (.A(_00432_),
    .B(_06599_),
    .ZN(_06774_));
 XNOR2_X1 _15947_ (.A(net539),
    .B(_06774_),
    .ZN(_06775_));
 OAI21_X1 _15948_ (.A(_06773_),
    .B1(_06775_),
    .B2(_06772_),
    .ZN(_00369_));
 BUF_X4 _15949_ (.A(_06771_),
    .Z(_06776_));
 NAND2_X1 _15950_ (.A1(_06776_),
    .A2(net150),
    .ZN(_06777_));
 XNOR2_X2 _15951_ (.A(_00433_),
    .B(_06615_),
    .ZN(_06778_));
 XNOR2_X1 _15952_ (.A(_06623_),
    .B(_06778_),
    .ZN(_06779_));
 OAI21_X1 _15953_ (.A(_06777_),
    .B1(_06779_),
    .B2(_06772_),
    .ZN(_00370_));
 NAND2_X1 _15954_ (.A1(_06776_),
    .A2(net151),
    .ZN(_06780_));
 XNOR2_X2 _15955_ (.A(_00434_),
    .B(_06631_),
    .ZN(_06781_));
 XNOR2_X1 _15956_ (.A(_06639_),
    .B(_06781_),
    .ZN(_06782_));
 OAI21_X1 _15957_ (.A(_06780_),
    .B1(_06782_),
    .B2(_06772_),
    .ZN(_00371_));
 NAND2_X1 _15958_ (.A1(_06776_),
    .A2(net158),
    .ZN(_06783_));
 XNOR2_X2 _15959_ (.A(_00435_),
    .B(_06652_),
    .ZN(_06784_));
 XNOR2_X1 _15960_ (.A(_06658_),
    .B(_06784_),
    .ZN(_06785_));
 OAI21_X1 _15961_ (.A(_06783_),
    .B1(_06785_),
    .B2(_06772_),
    .ZN(_00372_));
 NAND2_X1 _15962_ (.A1(_06776_),
    .A2(net164),
    .ZN(_06786_));
 XNOR2_X2 _15963_ (.A(_00436_),
    .B(_06667_),
    .ZN(_06787_));
 XNOR2_X1 _15964_ (.A(_06674_),
    .B(_06787_),
    .ZN(_06788_));
 OAI21_X1 _15965_ (.A(_06786_),
    .B1(_06788_),
    .B2(_06772_),
    .ZN(_00373_));
 NAND2_X1 _15966_ (.A1(_06776_),
    .A2(net167),
    .ZN(_06789_));
 XOR2_X2 _15967_ (.A(_00437_),
    .B(_06684_),
    .Z(_06790_));
 XNOR2_X1 _15968_ (.A(_06689_),
    .B(_06790_),
    .ZN(_06791_));
 OAI21_X1 _15969_ (.A(_06789_),
    .B1(_06791_),
    .B2(_06772_),
    .ZN(_00374_));
 XNOR2_X2 _15970_ (.A(_00438_),
    .B(_06702_),
    .ZN(_06792_));
 XNOR2_X1 _15971_ (.A(_06698_),
    .B(_06792_),
    .ZN(_06793_));
 MUX2_X1 _15972_ (.A(net168),
    .B(_06793_),
    .S(_06768_),
    .Z(_00376_));
 XNOR2_X2 _15973_ (.A(_00439_),
    .B(_06707_),
    .ZN(_06794_));
 XNOR2_X1 _15974_ (.A(_06711_),
    .B(_06794_),
    .ZN(_06795_));
 XOR2_X1 _15975_ (.A(_06710_),
    .B(_06795_),
    .Z(_06796_));
 MUX2_X1 _15976_ (.A(net169),
    .B(_06796_),
    .S(_06768_),
    .Z(_00377_));
 BUF_X4 _15977_ (.A(_06720_),
    .Z(_06797_));
 NOR2_X1 _15978_ (.A1(_06797_),
    .A2(net170),
    .ZN(_06798_));
 BUF_X4 _15979_ (.A(_06720_),
    .Z(_06799_));
 BUF_X4 _15980_ (.A(_06799_),
    .Z(_06800_));
 AOI21_X1 _15981_ (.A(_06798_),
    .B1(_06718_),
    .B2(_06800_),
    .ZN(_00321_));
 NOR2_X1 _15982_ (.A1(_06797_),
    .A2(net172),
    .ZN(_06801_));
 AOI21_X1 _15983_ (.A(_06801_),
    .B1(_06722_),
    .B2(_06800_),
    .ZN(_00332_));
 NOR2_X1 _15984_ (.A1(_06797_),
    .A2(net179),
    .ZN(_06802_));
 AOI21_X1 _15985_ (.A(_06802_),
    .B1(_06724_),
    .B2(_06800_),
    .ZN(_00343_));
 NOR2_X1 _15986_ (.A1(_06797_),
    .A2(net180),
    .ZN(_06803_));
 AOI21_X1 _15987_ (.A(_06803_),
    .B1(_06727_),
    .B2(_06800_),
    .ZN(_00346_));
 NOR2_X1 _15988_ (.A1(_06797_),
    .A2(net181),
    .ZN(_06804_));
 AOI21_X1 _15989_ (.A(_06804_),
    .B1(_06729_),
    .B2(_06800_),
    .ZN(_00347_));
 BUF_X4 _15990_ (.A(_06720_),
    .Z(_06805_));
 NOR2_X1 _15991_ (.A1(_06805_),
    .A2(net182),
    .ZN(_06806_));
 AOI21_X1 _15992_ (.A(_06806_),
    .B1(_06731_),
    .B2(_06800_),
    .ZN(_00348_));
 NOR2_X1 _15993_ (.A1(_06805_),
    .A2(net184),
    .ZN(_06807_));
 AOI21_X1 _15994_ (.A(_06807_),
    .B1(_06733_),
    .B2(_06800_),
    .ZN(_00349_));
 NOR2_X1 _15995_ (.A1(_06805_),
    .A2(net185),
    .ZN(_06808_));
 AOI21_X1 _15996_ (.A(_06808_),
    .B1(_06735_),
    .B2(_06800_),
    .ZN(_00350_));
 NOR2_X1 _15997_ (.A1(_06805_),
    .A2(net186),
    .ZN(_06809_));
 AOI21_X1 _15998_ (.A(_06809_),
    .B1(_06737_),
    .B2(_06800_),
    .ZN(_00351_));
 NOR2_X1 _15999_ (.A1(_06805_),
    .A2(net190),
    .ZN(_06810_));
 AOI21_X1 _16000_ (.A(_06810_),
    .B1(_06739_),
    .B2(_06800_),
    .ZN(_00352_));
 NOR2_X1 _16001_ (.A1(_06805_),
    .A2(net191),
    .ZN(_06811_));
 BUF_X4 _16002_ (.A(_06799_),
    .Z(_06812_));
 AOI21_X1 _16003_ (.A(_06811_),
    .B1(_06741_),
    .B2(_06812_),
    .ZN(_00322_));
 NOR2_X1 _16004_ (.A1(_06805_),
    .A2(net192),
    .ZN(_06813_));
 AOI21_X1 _16005_ (.A(_06813_),
    .B1(_06743_),
    .B2(_06812_),
    .ZN(_00323_));
 NOR2_X1 _16006_ (.A1(_06805_),
    .A2(net193),
    .ZN(_06814_));
 AOI21_X1 _16007_ (.A(_06814_),
    .B1(_06745_),
    .B2(_06812_),
    .ZN(_00324_));
 NOR2_X1 _16008_ (.A1(_06805_),
    .A2(net194),
    .ZN(_06815_));
 AOI21_X1 _16009_ (.A(_06815_),
    .B1(_06748_),
    .B2(_06812_),
    .ZN(_00325_));
 NOR2_X1 _16010_ (.A1(_06805_),
    .A2(net198),
    .ZN(_06816_));
 AOI21_X1 _16011_ (.A(_06816_),
    .B1(_06750_),
    .B2(_06812_),
    .ZN(_00326_));
 CLKBUF_X3 _16012_ (.A(_06720_),
    .Z(_06817_));
 NOR2_X1 _16013_ (.A1(_06817_),
    .A2(net199),
    .ZN(_06818_));
 AOI21_X1 _16014_ (.A(_06818_),
    .B1(_06752_),
    .B2(_06812_),
    .ZN(_00327_));
 NOR2_X1 _16015_ (.A1(_06817_),
    .A2(net204),
    .ZN(_06819_));
 AOI21_X1 _16016_ (.A(_06819_),
    .B1(_06754_),
    .B2(_06812_),
    .ZN(_00328_));
 NOR2_X1 _16017_ (.A1(_06817_),
    .A2(net205),
    .ZN(_06820_));
 AOI21_X1 _16018_ (.A(_06820_),
    .B1(_06756_),
    .B2(_06812_),
    .ZN(_00329_));
 MUX2_X1 _16019_ (.A(net206),
    .B(_06758_),
    .S(_06768_),
    .Z(_00330_));
 NOR2_X1 _16020_ (.A1(_06817_),
    .A2(net207),
    .ZN(_06821_));
 AOI21_X1 _16021_ (.A(_06821_),
    .B1(_06760_),
    .B2(_06812_),
    .ZN(_00331_));
 NOR2_X1 _16022_ (.A1(_06817_),
    .A2(net208),
    .ZN(_06822_));
 AOI21_X1 _16023_ (.A(_06822_),
    .B1(_06762_),
    .B2(_06812_),
    .ZN(_00333_));
 NOR2_X1 _16024_ (.A1(_06817_),
    .A2(net209),
    .ZN(_06823_));
 CLKBUF_X3 _16025_ (.A(_06799_),
    .Z(_06824_));
 AOI21_X1 _16026_ (.A(_06823_),
    .B1(_06764_),
    .B2(_06824_),
    .ZN(_00334_));
 NOR2_X1 _16027_ (.A1(_06817_),
    .A2(net210),
    .ZN(_06825_));
 AOI21_X1 _16028_ (.A(_06825_),
    .B1(_06766_),
    .B2(_06824_),
    .ZN(_00335_));
 NOR2_X1 _16029_ (.A1(_06817_),
    .A2(net211),
    .ZN(_06826_));
 AOI21_X1 _16030_ (.A(_06826_),
    .B1(_06769_),
    .B2(_06824_),
    .ZN(_00336_));
 XNOR2_X1 _16031_ (.A(net785),
    .B(_06774_),
    .ZN(_06827_));
 MUX2_X1 _16032_ (.A(net212),
    .B(_06827_),
    .S(_06768_),
    .Z(_00337_));
 XNOR2_X1 _16033_ (.A(net1088),
    .B(_06778_),
    .ZN(_06828_));
 MUX2_X1 _16034_ (.A(net213),
    .B(_06828_),
    .S(_06768_),
    .Z(_00338_));
 XNOR2_X1 _16035_ (.A(_06638_),
    .B(_06781_),
    .ZN(_06829_));
 MUX2_X1 _16036_ (.A(net215),
    .B(_06829_),
    .S(_06768_),
    .Z(_00339_));
 XNOR2_X1 _16037_ (.A(_06657_),
    .B(_06784_),
    .ZN(_06830_));
 MUX2_X1 _16038_ (.A(net216),
    .B(_06830_),
    .S(_06768_),
    .Z(_00340_));
 XNOR2_X1 _16039_ (.A(_06673_),
    .B(_06787_),
    .ZN(_06831_));
 MUX2_X1 _16040_ (.A(net217),
    .B(_06831_),
    .S(_06768_),
    .Z(_00341_));
 XNOR2_X1 _16041_ (.A(_06688_),
    .B(_06790_),
    .ZN(_06832_));
 BUF_X4 _16042_ (.A(_06720_),
    .Z(_06833_));
 MUX2_X1 _16043_ (.A(net218),
    .B(_06832_),
    .S(_06833_),
    .Z(_00342_));
 XNOR2_X1 _16044_ (.A(_06697_),
    .B(_06792_),
    .ZN(_06834_));
 MUX2_X1 _16045_ (.A(net219),
    .B(_06834_),
    .S(_06833_),
    .Z(_00344_));
 MUX2_X1 _16046_ (.A(net220),
    .B(_06795_),
    .S(_06833_),
    .Z(_00345_));
 XOR2_X1 _16047_ (.A(_06325_),
    .B(\u0.subword[0] ),
    .Z(_06835_));
 MUX2_X1 _16048_ (.A(net221),
    .B(_06835_),
    .S(_06833_),
    .Z(_00289_));
 XOR2_X1 _16049_ (.A(_06340_),
    .B(net828),
    .Z(_06836_));
 MUX2_X1 _16050_ (.A(net222),
    .B(_06836_),
    .S(_06833_),
    .Z(_00300_));
 XOR2_X1 _16051_ (.A(_06355_),
    .B(\u0.subword[2] ),
    .Z(_06837_));
 MUX2_X1 _16052_ (.A(net223),
    .B(_06837_),
    .S(_06833_),
    .Z(_00311_));
 XOR2_X1 _16053_ (.A(_06386_),
    .B(\u0.subword[3] ),
    .Z(_06838_));
 MUX2_X1 _16054_ (.A(net224),
    .B(_06838_),
    .S(_06833_),
    .Z(_00314_));
 XOR2_X1 _16055_ (.A(_06403_),
    .B(\u0.subword[4] ),
    .Z(_06839_));
 MUX2_X1 _16056_ (.A(net20),
    .B(_06839_),
    .S(_06833_),
    .Z(_00315_));
 XOR2_X1 _16057_ (.A(_06417_),
    .B(\u0.subword[5] ),
    .Z(_06840_));
 MUX2_X1 _16058_ (.A(net21),
    .B(_06840_),
    .S(_06833_),
    .Z(_00316_));
 XOR2_X1 _16059_ (.A(_06431_),
    .B(\u0.subword[6] ),
    .Z(_06841_));
 MUX2_X1 _16060_ (.A(net22),
    .B(_06841_),
    .S(_06833_),
    .Z(_00317_));
 XOR2_X1 _16061_ (.A(_06439_),
    .B(\u0.subword[7] ),
    .Z(_06842_));
 BUF_X4 _16062_ (.A(_06720_),
    .Z(_06843_));
 MUX2_X1 _16063_ (.A(net23),
    .B(_06842_),
    .S(_06843_),
    .Z(_00318_));
 XOR2_X1 _16064_ (.A(_06450_),
    .B(\u0.subword[8] ),
    .Z(_06844_));
 MUX2_X1 _16065_ (.A(net24),
    .B(_06844_),
    .S(_06843_),
    .Z(_00319_));
 XOR2_X1 _16066_ (.A(_06465_),
    .B(net1050),
    .Z(_06845_));
 MUX2_X1 _16067_ (.A(net25),
    .B(_06845_),
    .S(_06843_),
    .Z(_00320_));
 XOR2_X1 _16068_ (.A(_06480_),
    .B(\u0.subword[10] ),
    .Z(_06846_));
 MUX2_X1 _16069_ (.A(net26),
    .B(_06846_),
    .S(_06843_),
    .Z(_00290_));
 XOR2_X1 _16070_ (.A(_06510_),
    .B(\u0.subword[11] ),
    .Z(_06847_));
 MUX2_X1 _16071_ (.A(net30),
    .B(_06847_),
    .S(_06843_),
    .Z(_00291_));
 XOR2_X1 _16072_ (.A(_06527_),
    .B(\u0.subword[12] ),
    .Z(_06848_));
 MUX2_X1 _16073_ (.A(net31),
    .B(_06848_),
    .S(_06843_),
    .Z(_00292_));
 XOR2_X1 _16074_ (.A(_06542_),
    .B(\u0.subword[13] ),
    .Z(_06849_));
 MUX2_X1 _16075_ (.A(net33),
    .B(_06849_),
    .S(_06843_),
    .Z(_00293_));
 XOR2_X1 _16076_ (.A(_06555_),
    .B(\u0.subword[14] ),
    .Z(_06850_));
 MUX2_X1 _16077_ (.A(net35),
    .B(_06850_),
    .S(_06843_),
    .Z(_00294_));
 XOR2_X1 _16078_ (.A(_06564_),
    .B(\u0.subword[15] ),
    .Z(_06851_));
 MUX2_X1 _16079_ (.A(net38),
    .B(_06851_),
    .S(_06843_),
    .Z(_00295_));
 XOR2_X1 _16080_ (.A(_06241_),
    .B(\u0.subword[16] ),
    .Z(_06852_));
 MUX2_X1 _16081_ (.A(net40),
    .B(_06852_),
    .S(_06843_),
    .Z(_00296_));
 XOR2_X1 _16082_ (.A(_06255_),
    .B(\u0.subword[17] ),
    .Z(_06853_));
 MUX2_X1 _16083_ (.A(net41),
    .B(_06853_),
    .S(_06799_),
    .Z(_00297_));
 XOR2_X1 _16084_ (.A(net1003),
    .B(\u0.subword[18] ),
    .Z(_06854_));
 MUX2_X1 _16085_ (.A(net44),
    .B(_06854_),
    .S(_06799_),
    .Z(_00298_));
 XOR2_X1 _16086_ (.A(_06221_),
    .B(\u0.subword[19] ),
    .Z(_06855_));
 MUX2_X1 _16087_ (.A(net45),
    .B(_06855_),
    .S(_06799_),
    .Z(_00299_));
 XOR2_X1 _16088_ (.A(_06281_),
    .B(\u0.subword[20] ),
    .Z(_06856_));
 MUX2_X1 _16089_ (.A(net46),
    .B(_06856_),
    .S(_06799_),
    .Z(_00301_));
 XOR2_X1 _16090_ (.A(_06269_),
    .B(\u0.subword[21] ),
    .Z(_06857_));
 MUX2_X1 _16091_ (.A(net47),
    .B(_06857_),
    .S(_06799_),
    .Z(_00302_));
 XOR2_X1 _16092_ (.A(_06575_),
    .B(\u0.subword[22] ),
    .Z(_06858_));
 MUX2_X1 _16093_ (.A(net48),
    .B(_06858_),
    .S(_06799_),
    .Z(_00303_));
 XOR2_X1 _16094_ (.A(_06587_),
    .B(\u0.subword[23] ),
    .Z(_06859_));
 MUX2_X1 _16095_ (.A(net50),
    .B(_06859_),
    .S(_06799_),
    .Z(_00304_));
 NOR2_X1 _16096_ (.A1(_06817_),
    .A2(net53),
    .ZN(_06860_));
 AOI21_X1 _16097_ (.A(_06860_),
    .B1(_06774_),
    .B2(_06824_),
    .ZN(_00305_));
 NOR2_X1 _16098_ (.A1(_06817_),
    .A2(net54),
    .ZN(_06861_));
 AOI21_X1 _16099_ (.A(_06861_),
    .B1(_06778_),
    .B2(_06824_),
    .ZN(_00306_));
 NOR2_X1 _16100_ (.A1(_06721_),
    .A2(net55),
    .ZN(_06862_));
 AOI21_X1 _16101_ (.A(_06862_),
    .B1(_06781_),
    .B2(_06824_),
    .ZN(_00307_));
 NOR2_X1 _16102_ (.A1(_06721_),
    .A2(net56),
    .ZN(_06863_));
 AOI21_X1 _16103_ (.A(_06863_),
    .B1(_06784_),
    .B2(_06824_),
    .ZN(_00308_));
 NOR2_X1 _16104_ (.A1(_06721_),
    .A2(net58),
    .ZN(_06864_));
 AOI21_X2 _16105_ (.A(_06864_),
    .B1(_06787_),
    .B2(_06824_),
    .ZN(_00309_));
 NOR2_X1 _16106_ (.A1(_06721_),
    .A2(net59),
    .ZN(_06865_));
 AOI21_X1 _16107_ (.A(_06865_),
    .B1(_06790_),
    .B2(_06824_),
    .ZN(_00310_));
 NOR2_X1 _16108_ (.A1(_06721_),
    .A2(net60),
    .ZN(_06866_));
 AOI21_X1 _16109_ (.A(_06866_),
    .B1(_06792_),
    .B2(_06824_),
    .ZN(_00312_));
 NOR2_X1 _16110_ (.A1(_06721_),
    .A2(net61),
    .ZN(_06867_));
 AOI21_X2 _16111_ (.A(_06867_),
    .B1(_06794_),
    .B2(_06797_),
    .ZN(_00313_));
 BUF_X8 _16112_ (.A(_06265_),
    .Z(_06868_));
 BUF_X2 clone361 (.A(net879),
    .Z(net878));
 BUF_X16 _16114_ (.A(_06319_),
    .Z(_06869_));
 BUF_X8 _16115_ (.A(_06869_),
    .Z(_06870_));
 BUF_X4 rebuffer470 (.A(_15306_),
    .Z(net1028));
 BUF_X16 _16117_ (.A(_06870_),
    .Z(_14678_));
 BUF_X8 _16118_ (.A(_06252_),
    .Z(_14659_));
 NOR2_X1 _16119_ (.A1(_06277_),
    .A2(_06596_),
    .ZN(_06872_));
 BUF_X4 _16120_ (.A(_06583_),
    .Z(_06873_));
 CLKBUF_X3 _16121_ (.A(_06873_),
    .Z(_06874_));
 NOR2_X2 clone42 (.A1(_06264_),
    .A2(_06254_),
    .ZN(net42));
 INV_X2 _16123_ (.A(_14661_),
    .ZN(_06876_));
 NAND2_X2 _16124_ (.A1(net43),
    .A2(_06323_),
    .ZN(_06877_));
 CLKBUF_X2 _16125_ (.A(_14660_),
    .Z(_06878_));
 CLKBUF_X3 _16126_ (.A(_06878_),
    .Z(_06879_));
 BUF_X8 _16127_ (.A(net999),
    .Z(_06880_));
 BUF_X4 _16128_ (.A(_06880_),
    .Z(_06881_));
 NAND2_X1 _16129_ (.A1(_06879_),
    .A2(_06881_),
    .ZN(_06882_));
 BUF_X4 _16130_ (.A(_06236_),
    .Z(_06883_));
 NOR2_X1 _16131_ (.A1(_06883_),
    .A2(_06291_),
    .ZN(_06884_));
 NAND3_X1 _16132_ (.A1(_06877_),
    .A2(_06882_),
    .A3(_06884_),
    .ZN(_06885_));
 BUF_X4 _16133_ (.A(_06233_),
    .Z(_06886_));
 NOR2_X4 _16134_ (.A1(_06886_),
    .A2(_06291_),
    .ZN(_06887_));
 BUF_X1 rebuffer741 (.A(_14661_),
    .Z(net1204));
 NAND2_X1 _16136_ (.A1(_14674_),
    .A2(_06880_),
    .ZN(_06889_));
 BUF_X4 _16137_ (.A(_14670_),
    .Z(_06890_));
 NAND2_X1 _16138_ (.A1(_06890_),
    .A2(_06322_),
    .ZN(_06891_));
 NAND3_X1 _16139_ (.A1(_06887_),
    .A2(_06889_),
    .A3(_06891_),
    .ZN(_06892_));
 NAND3_X1 _16140_ (.A1(_06874_),
    .A2(_06885_),
    .A3(_06892_),
    .ZN(_06893_));
 OAI22_X4 _16141_ (.A1(_06240_),
    .A2(_06251_),
    .B1(_06254_),
    .B2(_06264_),
    .ZN(_06894_));
 OAI211_X2 _16142_ (.A(_06883_),
    .B(_06894_),
    .C1(_06881_),
    .C2(_14664_),
    .ZN(_06895_));
 BUF_X4 _16143_ (.A(_06233_),
    .Z(_06896_));
 BUF_X4 _16144_ (.A(_06896_),
    .Z(_06897_));
 CLKBUF_X3 _16145_ (.A(_06897_),
    .Z(_06898_));
 NOR2_X2 _16146_ (.A1(net801),
    .A2(net64),
    .ZN(_06899_));
 NOR2_X1 _16147_ (.A1(net1000),
    .A2(_06881_),
    .ZN(_06900_));
 OAI21_X1 _16148_ (.A(_06898_),
    .B1(_06899_),
    .B2(_06900_),
    .ZN(_06901_));
 AND3_X1 _16149_ (.A1(_00391_),
    .A2(_06895_),
    .A3(_06901_),
    .ZN(_06902_));
 BUF_X4 _16150_ (.A(_06289_),
    .Z(_06903_));
 BUF_X4 _16151_ (.A(_06903_),
    .Z(_06904_));
 CLKBUF_X3 _16152_ (.A(_06904_),
    .Z(_06905_));
 BUF_X4 clone64 (.A(net615),
    .Z(net64));
 INV_X2 _16154_ (.A(_14665_),
    .ZN(_06907_));
 NOR2_X1 _16155_ (.A1(net65),
    .A2(_14683_),
    .ZN(_06908_));
 BUF_X4 clone94 (.A(net1158),
    .Z(net94));
 CLKBUF_X3 _16157_ (.A(_14667_),
    .Z(_06910_));
 NOR2_X2 _16158_ (.A1(_06910_),
    .A2(_06881_),
    .ZN(_06911_));
 OAI21_X1 _16159_ (.A(_00390_),
    .B1(_06908_),
    .B2(_06911_),
    .ZN(_06912_));
 NAND2_X2 _16160_ (.A1(net1000),
    .A2(_06870_),
    .ZN(_06913_));
 OAI21_X1 _16161_ (.A(_06912_),
    .B1(_06913_),
    .B2(_00390_),
    .ZN(_06914_));
 BUF_X4 _16162_ (.A(net1194),
    .Z(_06915_));
 BUF_X4 _16163_ (.A(_06319_),
    .Z(_06916_));
 BUF_X4 _16164_ (.A(_06916_),
    .Z(_06917_));
 NAND2_X2 _16165_ (.A1(_06915_),
    .A2(_06917_),
    .ZN(_06918_));
 CLKBUF_X3 _16166_ (.A(_06235_),
    .Z(_06919_));
 NOR2_X4 _16167_ (.A1(net518),
    .A2(_06319_),
    .ZN(_06920_));
 NOR2_X2 _16168_ (.A1(_06919_),
    .A2(_06920_),
    .ZN(_06921_));
 AOI21_X2 _16169_ (.A(_06905_),
    .B1(_06918_),
    .B2(_06921_),
    .ZN(_06922_));
 BUF_X4 rebuffer406 (.A(\sa12_sr[1] ),
    .Z(net930));
 INV_X2 _16171_ (.A(_14662_),
    .ZN(_06924_));
 NAND2_X2 _16172_ (.A1(_06924_),
    .A2(_06916_),
    .ZN(_06925_));
 NAND3_X1 _16173_ (.A1(_00390_),
    .A2(_06877_),
    .A3(_06925_),
    .ZN(_06926_));
 AOI22_X2 _16174_ (.A1(_06905_),
    .A2(_06914_),
    .B1(_06922_),
    .B2(_06926_),
    .ZN(_06927_));
 OAI221_X2 _16175_ (.A(_06872_),
    .B1(_06893_),
    .B2(_06902_),
    .C1(_06927_),
    .C2(_06874_),
    .ZN(_06928_));
 BUF_X4 _16176_ (.A(_06595_),
    .Z(_06929_));
 NOR2_X2 _16177_ (.A1(_06277_),
    .A2(_06929_),
    .ZN(_06930_));
 BUF_X8 _16178_ (.A(_06321_),
    .Z(_06931_));
 BUF_X4 _16179_ (.A(_06931_),
    .Z(_06932_));
 NAND2_X1 _16180_ (.A1(_06915_),
    .A2(_06932_),
    .ZN(_06933_));
 CLKBUF_X3 _16181_ (.A(_14672_),
    .Z(_06934_));
 INV_X2 _16182_ (.A(_06934_),
    .ZN(_06935_));
 NAND2_X1 _16183_ (.A1(_06935_),
    .A2(_14678_),
    .ZN(_06936_));
 NAND3_X1 _16184_ (.A1(_06887_),
    .A2(_06933_),
    .A3(_06936_),
    .ZN(_06937_));
 NAND2_X2 _16185_ (.A1(_06233_),
    .A2(_06290_),
    .ZN(_06938_));
 BUF_X1 rebuffer730 (.A(_14665_),
    .Z(net1193));
 NAND2_X1 _16187_ (.A1(net1195),
    .A2(_14683_),
    .ZN(_06940_));
 NOR2_X1 _16188_ (.A1(_06887_),
    .A2(_06940_),
    .ZN(_06941_));
 NOR2_X2 _16189_ (.A1(_06883_),
    .A2(_06903_),
    .ZN(_06942_));
 NAND2_X2 _16190_ (.A1(_06890_),
    .A2(_06916_),
    .ZN(_06943_));
 AND2_X1 _16191_ (.A1(_06942_),
    .A2(_06943_),
    .ZN(_06944_));
 AOI22_X1 _16192_ (.A1(_06938_),
    .A2(_06941_),
    .B1(_06933_),
    .B2(_06944_),
    .ZN(_06945_));
 NAND3_X1 _16193_ (.A1(_06874_),
    .A2(_06937_),
    .A3(_06945_),
    .ZN(_06946_));
 NAND2_X1 _16194_ (.A1(_06930_),
    .A2(_06946_),
    .ZN(_06947_));
 CLKBUF_X3 _16195_ (.A(_06919_),
    .Z(_06948_));
 CLKBUF_X3 _16196_ (.A(_06948_),
    .Z(_06949_));
 MUX2_X1 _16197_ (.A(_14661_),
    .B(_06265_),
    .S(_06321_),
    .Z(_06950_));
 NOR2_X1 _16198_ (.A1(_06949_),
    .A2(_06950_),
    .ZN(_06951_));
 CLKBUF_X3 _16199_ (.A(_06886_),
    .Z(_06952_));
 CLKBUF_X3 _16200_ (.A(_06952_),
    .Z(_06953_));
 NAND2_X2 _16201_ (.A1(net802),
    .A2(_06931_),
    .ZN(_06954_));
 INV_X1 _16202_ (.A(_06890_),
    .ZN(_06955_));
 NAND2_X1 _16203_ (.A1(_06955_),
    .A2(_06870_),
    .ZN(_06956_));
 AOI21_X1 _16204_ (.A(_06953_),
    .B1(_06954_),
    .B2(_06956_),
    .ZN(_06957_));
 NOR3_X1 _16205_ (.A1(_00391_),
    .A2(_06951_),
    .A3(_06957_),
    .ZN(_06958_));
 INV_X1 _16206_ (.A(_14674_),
    .ZN(_06959_));
 MUX2_X1 _16207_ (.A(net1195),
    .B(_06959_),
    .S(_06870_),
    .Z(_06960_));
 NAND2_X1 _16208_ (.A1(_06236_),
    .A2(_06932_),
    .ZN(_06961_));
 OAI22_X1 _16209_ (.A1(_00390_),
    .A2(_06960_),
    .B1(_06961_),
    .B2(_06910_),
    .ZN(_06962_));
 AOI21_X1 _16210_ (.A(_06958_),
    .B1(_06962_),
    .B2(_00391_),
    .ZN(_06963_));
 NOR2_X1 _16211_ (.A1(_06874_),
    .A2(_06963_),
    .ZN(_06964_));
 CLKBUF_X3 _16212_ (.A(net517),
    .Z(_06965_));
 MUX2_X1 _16213_ (.A(_06915_),
    .B(_06965_),
    .S(_06880_),
    .Z(_06966_));
 MUX2_X1 _16214_ (.A(_14674_),
    .B(_06253_),
    .S(_06880_),
    .Z(_06967_));
 MUX2_X1 _16215_ (.A(_06966_),
    .B(_06967_),
    .S(_06883_),
    .Z(_06968_));
 INV_X1 _16216_ (.A(_14667_),
    .ZN(_06969_));
 NOR2_X2 _16217_ (.A1(_06969_),
    .A2(_06235_),
    .ZN(_06970_));
 INV_X2 _16218_ (.A(_06878_),
    .ZN(_06971_));
 MUX2_X1 _16219_ (.A(_06971_),
    .B(_06965_),
    .S(_06880_),
    .Z(_06972_));
 AOI221_X2 _16220_ (.A(_06292_),
    .B1(_06881_),
    .B2(_06970_),
    .C1(_06972_),
    .C2(_06237_),
    .ZN(_06973_));
 MUX2_X1 _16221_ (.A(_06968_),
    .B(_06973_),
    .S(_06585_),
    .Z(_06974_));
 NOR2_X1 _16222_ (.A1(_00391_),
    .A2(_06974_),
    .ZN(_06975_));
 MUX2_X1 _16223_ (.A(_06910_),
    .B(_06934_),
    .S(_06323_),
    .Z(_06976_));
 NOR2_X1 _16224_ (.A1(_06949_),
    .A2(_06976_),
    .ZN(_06977_));
 BUF_X2 _16225_ (.A(_14661_),
    .Z(_06978_));
 NOR3_X2 _16226_ (.A1(net51),
    .A2(_06896_),
    .A3(_06917_),
    .ZN(_06979_));
 NOR4_X2 _16227_ (.A1(_06874_),
    .A2(_06973_),
    .A3(_06977_),
    .A4(_06979_),
    .ZN(_06980_));
 OAI21_X1 _16228_ (.A(_06873_),
    .B1(_06897_),
    .B2(_14686_),
    .ZN(_06981_));
 NAND2_X2 _16229_ (.A1(_06978_),
    .A2(_06881_),
    .ZN(_06982_));
 AOI221_X2 _16230_ (.A(_06981_),
    .B1(_06968_),
    .B2(_06904_),
    .C1(_06898_),
    .C2(_06982_),
    .ZN(_06983_));
 NOR4_X2 _16231_ (.A1(_06929_),
    .A2(_06975_),
    .A3(_06980_),
    .A4(_06983_),
    .ZN(_06984_));
 BUF_X4 _16232_ (.A(_06277_),
    .Z(_06985_));
 BUF_X4 _16233_ (.A(_06903_),
    .Z(_06986_));
 MUX2_X1 _16234_ (.A(_06878_),
    .B(_14664_),
    .S(_06870_),
    .Z(_06987_));
 OAI21_X1 _16235_ (.A(_06986_),
    .B1(_06987_),
    .B2(_06952_),
    .ZN(_06988_));
 NAND2_X2 _16236_ (.A1(_14669_),
    .A2(_06917_),
    .ZN(_06989_));
 AOI21_X1 _16237_ (.A(_06238_),
    .B1(_06940_),
    .B2(_06989_),
    .ZN(_06990_));
 MUX2_X1 _16238_ (.A(net65),
    .B(_06868_),
    .S(_06322_),
    .Z(_06991_));
 MUX2_X1 _16239_ (.A(_14662_),
    .B(_14659_),
    .S(_06870_),
    .Z(_06992_));
 MUX2_X1 _16240_ (.A(_06991_),
    .B(_06992_),
    .S(_06238_),
    .Z(_06993_));
 OAI221_X1 _16241_ (.A(_00393_),
    .B1(_06988_),
    .B2(_06990_),
    .C1(_06993_),
    .C2(_06905_),
    .ZN(_06994_));
 CLKBUF_X3 _16242_ (.A(_06292_),
    .Z(_06995_));
 BUF_X4 _16243_ (.A(_06995_),
    .Z(_06996_));
 NOR2_X1 _16244_ (.A1(_06868_),
    .A2(_06931_),
    .ZN(_06997_));
 BUF_X8 _16245_ (.A(_06978_),
    .Z(_06998_));
 NAND2_X1 _16246_ (.A1(_06998_),
    .A2(_06953_),
    .ZN(_06999_));
 OAI21_X1 _16247_ (.A(_14678_),
    .B1(net66),
    .B2(_06238_),
    .ZN(_07000_));
 OAI221_X1 _16248_ (.A(_06996_),
    .B1(_06997_),
    .B2(_06999_),
    .C1(_07000_),
    .C2(_06998_),
    .ZN(_07001_));
 NOR2_X4 _16249_ (.A1(_06235_),
    .A2(_06931_),
    .ZN(_07002_));
 XNOR2_X2 _16250_ (.A(_06234_),
    .B(net999),
    .ZN(_07003_));
 CLKBUF_X3 _16251_ (.A(_14674_),
    .Z(_07004_));
 AOI221_X1 _16252_ (.A(_06979_),
    .B1(_07002_),
    .B2(_06890_),
    .C1(_07003_),
    .C2(_07004_),
    .ZN(_07005_));
 OAI21_X1 _16253_ (.A(_07001_),
    .B1(_07005_),
    .B2(_00391_),
    .ZN(_07006_));
 OAI21_X1 _16254_ (.A(_06994_),
    .B1(_07006_),
    .B2(_00393_),
    .ZN(_07007_));
 OAI21_X1 _16255_ (.A(_06985_),
    .B1(_00394_),
    .B2(_07007_),
    .ZN(_07008_));
 OAI221_X2 _16256_ (.A(_06928_),
    .B1(_06947_),
    .B2(_06964_),
    .C1(_06984_),
    .C2(_07008_),
    .ZN(_00000_));
 MUX2_X1 _16257_ (.A(_14674_),
    .B(_06253_),
    .S(_06931_),
    .Z(_07009_));
 MUX2_X1 _16258_ (.A(_06878_),
    .B(net1194),
    .S(_06880_),
    .Z(_07010_));
 MUX2_X1 _16259_ (.A(_07009_),
    .B(_07010_),
    .S(_06883_),
    .Z(_07011_));
 MUX2_X1 _16260_ (.A(_06969_),
    .B(_14669_),
    .S(_06916_),
    .Z(_07012_));
 MUX2_X1 _16261_ (.A(_06965_),
    .B(net42),
    .S(_06880_),
    .Z(_07013_));
 MUX2_X1 _16262_ (.A(_07012_),
    .B(_07013_),
    .S(_06896_),
    .Z(_07014_));
 MUX2_X1 _16263_ (.A(_07011_),
    .B(_07014_),
    .S(_06277_),
    .Z(_07015_));
 OAI21_X1 _16264_ (.A(_06943_),
    .B1(_06870_),
    .B2(_06971_),
    .ZN(_07016_));
 OR2_X1 _16265_ (.A1(_14688_),
    .A2(_06278_),
    .ZN(_07017_));
 CLKBUF_X3 _16266_ (.A(_06237_),
    .Z(_07018_));
 MUX2_X1 _16267_ (.A(_07016_),
    .B(_07017_),
    .S(_07018_),
    .Z(_07019_));
 MUX2_X1 _16268_ (.A(_07015_),
    .B(_07019_),
    .S(_06904_),
    .Z(_07020_));
 OAI21_X2 _16269_ (.A(_06894_),
    .B1(net999),
    .B2(_14669_),
    .ZN(_07021_));
 NAND2_X2 _16270_ (.A1(_06883_),
    .A2(_06881_),
    .ZN(_07022_));
 OAI221_X1 _16271_ (.A(_06904_),
    .B1(_07021_),
    .B2(_06948_),
    .C1(_07022_),
    .C2(_06915_),
    .ZN(_07023_));
 MUX2_X1 _16272_ (.A(_06978_),
    .B(_06965_),
    .S(_06870_),
    .Z(_07024_));
 MUX2_X1 _16273_ (.A(_06910_),
    .B(_14664_),
    .S(_06917_),
    .Z(_07025_));
 MUX2_X1 _16274_ (.A(_07024_),
    .B(_07025_),
    .S(_06952_),
    .Z(_07026_));
 OAI21_X1 _16275_ (.A(_07023_),
    .B1(_07026_),
    .B2(_06904_),
    .ZN(_07027_));
 OAI21_X1 _16276_ (.A(_06886_),
    .B1(_06322_),
    .B2(_14667_),
    .ZN(_07028_));
 MUX2_X1 _16277_ (.A(net1193),
    .B(_06265_),
    .S(_06290_),
    .Z(_07029_));
 AOI21_X1 _16278_ (.A(_07028_),
    .B1(_07029_),
    .B2(_06932_),
    .ZN(_07030_));
 NOR2_X1 _16279_ (.A1(_14679_),
    .A2(_06903_),
    .ZN(_07031_));
 NAND2_X2 _16280_ (.A1(_14669_),
    .A2(_06931_),
    .ZN(_07032_));
 AOI21_X1 _16281_ (.A(_06235_),
    .B1(_06870_),
    .B2(_06910_),
    .ZN(_07033_));
 NAND2_X1 _16282_ (.A1(_07032_),
    .A2(_07033_),
    .ZN(_07034_));
 MUX2_X1 _16283_ (.A(net51),
    .B(_14662_),
    .S(_06322_),
    .Z(_07035_));
 AOI221_X1 _16284_ (.A(_07030_),
    .B1(_07031_),
    .B2(_07034_),
    .C1(_06887_),
    .C2(_07035_),
    .ZN(_07036_));
 MUX2_X1 _16285_ (.A(_07027_),
    .B(_07036_),
    .S(_06985_),
    .Z(_07037_));
 MUX2_X1 _16286_ (.A(_07020_),
    .B(_07037_),
    .S(_00394_),
    .Z(_07038_));
 NAND2_X1 _16287_ (.A1(_06924_),
    .A2(_14683_),
    .ZN(_07039_));
 OAI221_X1 _16288_ (.A(_07039_),
    .B1(_06232_),
    .B2(_06219_),
    .C1(net1195),
    .C2(_14683_),
    .ZN(_07040_));
 NAND2_X2 _16289_ (.A1(_06998_),
    .A2(_06932_),
    .ZN(_07041_));
 NAND3_X1 _16290_ (.A1(_06949_),
    .A2(_07041_),
    .A3(_06882_),
    .ZN(_07042_));
 AND3_X1 _16291_ (.A1(_06996_),
    .A2(_07040_),
    .A3(_07042_),
    .ZN(_07043_));
 AOI21_X1 _16292_ (.A(_06979_),
    .B1(_06987_),
    .B2(_06898_),
    .ZN(_07044_));
 NOR2_X1 _16293_ (.A1(_00391_),
    .A2(_07044_),
    .ZN(_07045_));
 NOR3_X1 _16294_ (.A1(_00392_),
    .A2(_07043_),
    .A3(_07045_),
    .ZN(_07046_));
 OAI221_X1 _16295_ (.A(_06913_),
    .B1(_06232_),
    .B2(_06219_),
    .C1(net1196),
    .C2(_14678_),
    .ZN(_07047_));
 NAND2_X2 _16296_ (.A1(_06876_),
    .A2(_06880_),
    .ZN(_07048_));
 NAND2_X1 _16297_ (.A1(_07004_),
    .A2(_06323_),
    .ZN(_07049_));
 NAND3_X1 _16298_ (.A1(_06949_),
    .A2(_07048_),
    .A3(_07049_),
    .ZN(_07050_));
 NAND3_X1 _16299_ (.A1(_00391_),
    .A2(_07047_),
    .A3(_07050_),
    .ZN(_07051_));
 AND2_X1 _16300_ (.A1(_06949_),
    .A2(_07012_),
    .ZN(_07052_));
 NOR2_X1 _16301_ (.A1(_07004_),
    .A2(_14683_),
    .ZN(_07053_));
 NOR3_X1 _16302_ (.A1(_06949_),
    .A2(_06920_),
    .A3(_07053_),
    .ZN(_07054_));
 OAI21_X1 _16303_ (.A(_06904_),
    .B1(_07052_),
    .B2(_07054_),
    .ZN(_07055_));
 AND3_X1 _16304_ (.A1(_00392_),
    .A2(_07051_),
    .A3(_07055_),
    .ZN(_07056_));
 OAI21_X1 _16305_ (.A(_06929_),
    .B1(_07046_),
    .B2(_07056_),
    .ZN(_07057_));
 NAND2_X1 _16306_ (.A1(_06905_),
    .A2(_06930_),
    .ZN(_07058_));
 NAND3_X1 _16307_ (.A1(_06910_),
    .A2(_06898_),
    .A3(_14683_),
    .ZN(_07059_));
 AOI21_X1 _16308_ (.A(_07058_),
    .B1(_07059_),
    .B2(_07042_),
    .ZN(_07060_));
 MUX2_X1 _16309_ (.A(_06998_),
    .B(_06969_),
    .S(_06881_),
    .Z(_07061_));
 NOR2_X4 _16310_ (.A1(_06886_),
    .A2(_06289_),
    .ZN(_07062_));
 AOI22_X1 _16311_ (.A1(_06942_),
    .A2(_06967_),
    .B1(_07061_),
    .B2(_07062_),
    .ZN(_07063_));
 NAND3_X1 _16312_ (.A1(_06985_),
    .A2(_00394_),
    .A3(_07063_),
    .ZN(_07064_));
 NAND2_X1 _16313_ (.A1(net1000),
    .A2(_06322_),
    .ZN(_07065_));
 NAND3_X1 _16314_ (.A1(_06898_),
    .A2(_07065_),
    .A3(_06982_),
    .ZN(_07066_));
 NAND2_X1 _16315_ (.A1(_06965_),
    .A2(_14669_),
    .ZN(_07067_));
 NAND3_X1 _16316_ (.A1(_00390_),
    .A2(_06913_),
    .A3(_07067_),
    .ZN(_07068_));
 AOI21_X1 _16317_ (.A(_07064_),
    .B1(_07066_),
    .B2(_07068_),
    .ZN(_07069_));
 NAND2_X2 _16318_ (.A1(_06896_),
    .A2(_06932_),
    .ZN(_07070_));
 NOR2_X1 _16319_ (.A1(_06879_),
    .A2(_07070_),
    .ZN(_07071_));
 AND3_X1 _16320_ (.A1(_07018_),
    .A2(_06925_),
    .A3(_07032_),
    .ZN(_07072_));
 OAI21_X1 _16321_ (.A(_06930_),
    .B1(_07071_),
    .B2(_07072_),
    .ZN(_07073_));
 AOI21_X1 _16322_ (.A(_06905_),
    .B1(_07064_),
    .B2(_07073_),
    .ZN(_07074_));
 NOR4_X2 _16323_ (.A1(_07074_),
    .A2(_07060_),
    .A3(_07069_),
    .A4(_06874_),
    .ZN(_07075_));
 AOI22_X2 _16324_ (.A1(_07038_),
    .A2(_06874_),
    .B1(_07057_),
    .B2(_07075_),
    .ZN(_00001_));
 MUX2_X1 _16325_ (.A(_06907_),
    .B(_14669_),
    .S(_06321_),
    .Z(_07076_));
 MUX2_X1 _16326_ (.A(_14681_),
    .B(_07076_),
    .S(_06236_),
    .Z(_07077_));
 AOI22_X1 _16327_ (.A1(_14684_),
    .A2(_06237_),
    .B1(_07002_),
    .B2(_06915_),
    .ZN(_07078_));
 MUX2_X1 _16328_ (.A(_07077_),
    .B(_07078_),
    .S(_06986_),
    .Z(_07079_));
 NOR3_X1 _16329_ (.A1(_06890_),
    .A2(_06235_),
    .A3(_06931_),
    .ZN(_07080_));
 AOI221_X2 _16330_ (.A(_07080_),
    .B1(_06920_),
    .B2(_06236_),
    .C1(_06971_),
    .C2(_07003_),
    .ZN(_07081_));
 MUX2_X1 _16331_ (.A(net51),
    .B(_06910_),
    .S(_06917_),
    .Z(_07082_));
 NAND2_X1 _16332_ (.A1(_06948_),
    .A2(_07082_),
    .ZN(_07083_));
 NOR3_X1 _16333_ (.A1(_07004_),
    .A2(_06919_),
    .A3(_06917_),
    .ZN(_07084_));
 NOR2_X1 _16334_ (.A1(_06995_),
    .A2(_07084_),
    .ZN(_07085_));
 AOI22_X1 _16335_ (.A1(_06293_),
    .A2(_07081_),
    .B1(_07083_),
    .B2(_07085_),
    .ZN(_07086_));
 MUX2_X1 _16336_ (.A(_07079_),
    .B(_07086_),
    .S(_06278_),
    .Z(_07087_));
 MUX2_X1 _16337_ (.A(_14662_),
    .B(_14667_),
    .S(_06321_),
    .Z(_07088_));
 MUX2_X1 _16338_ (.A(_07076_),
    .B(_07088_),
    .S(_06886_),
    .Z(_07089_));
 MUX2_X1 _16339_ (.A(_14667_),
    .B(_06907_),
    .S(_06321_),
    .Z(_07090_));
 MUX2_X1 _16340_ (.A(_06950_),
    .B(_07090_),
    .S(_06236_),
    .Z(_07091_));
 MUX2_X1 _16341_ (.A(_07089_),
    .B(_07091_),
    .S(_06986_),
    .Z(_07092_));
 MUX2_X1 _16342_ (.A(net1204),
    .B(_14669_),
    .S(_06869_),
    .Z(_07093_));
 MUX2_X1 _16343_ (.A(_14676_),
    .B(_06252_),
    .S(_06321_),
    .Z(_07094_));
 MUX2_X1 _16344_ (.A(_07093_),
    .B(_07094_),
    .S(_06236_),
    .Z(_07095_));
 MUX2_X1 _16345_ (.A(_06924_),
    .B(_06878_),
    .S(_06916_),
    .Z(_07096_));
 AOI22_X1 _16346_ (.A1(_06915_),
    .A2(_07002_),
    .B1(_07096_),
    .B2(_06883_),
    .ZN(_07097_));
 MUX2_X1 _16347_ (.A(_07095_),
    .B(_07097_),
    .S(_06986_),
    .Z(_07098_));
 MUX2_X1 _16348_ (.A(_07092_),
    .B(_07098_),
    .S(_06278_),
    .Z(_07099_));
 MUX2_X1 _16349_ (.A(_07087_),
    .B(_07099_),
    .S(_06929_),
    .Z(_07100_));
 AOI21_X1 _16350_ (.A(_06938_),
    .B1(_06925_),
    .B2(_07065_),
    .ZN(_07101_));
 NAND2_X1 _16351_ (.A1(_06934_),
    .A2(_06323_),
    .ZN(_07102_));
 NAND3_X1 _16352_ (.A1(_07062_),
    .A2(_06989_),
    .A3(_07102_),
    .ZN(_07103_));
 NAND2_X1 _16353_ (.A1(_00392_),
    .A2(_07103_),
    .ZN(_07104_));
 XNOR2_X2 _16354_ (.A(net999),
    .B(_06876_),
    .ZN(_07105_));
 MUX2_X1 _16355_ (.A(_06934_),
    .B(_06965_),
    .S(_06322_),
    .Z(_07106_));
 MUX2_X1 _16356_ (.A(_07105_),
    .B(_07106_),
    .S(_06896_),
    .Z(_07107_));
 NOR2_X2 _16357_ (.A1(_06293_),
    .A2(_07107_),
    .ZN(_07108_));
 AOI21_X1 _16358_ (.A(_06938_),
    .B1(_06870_),
    .B2(_14662_),
    .ZN(_07109_));
 AND2_X1 _16359_ (.A1(_07102_),
    .A2(_07109_),
    .ZN(_07110_));
 AOI21_X1 _16360_ (.A(_06903_),
    .B1(_06954_),
    .B2(_06236_),
    .ZN(_07111_));
 NOR2_X4 _16361_ (.A1(_06290_),
    .A2(_06916_),
    .ZN(_07112_));
 MUX2_X1 _16362_ (.A(_06934_),
    .B(net42),
    .S(_06235_),
    .Z(_07113_));
 AOI221_X1 _16363_ (.A(_07111_),
    .B1(_07112_),
    .B2(_07113_),
    .C1(_06870_),
    .C2(_06910_),
    .ZN(_07114_));
 OAI33_X1 _16364_ (.A1(_07101_),
    .A2(_07104_),
    .A3(_07108_),
    .B1(_07110_),
    .B2(_07114_),
    .B3(_00392_),
    .ZN(_07115_));
 AOI21_X1 _16365_ (.A(_06938_),
    .B1(_07032_),
    .B2(_06889_),
    .ZN(_07116_));
 MUX2_X1 _16366_ (.A(_14688_),
    .B(_07021_),
    .S(_06235_),
    .Z(_07117_));
 NAND2_X1 _16367_ (.A1(_06891_),
    .A2(_07048_),
    .ZN(_07118_));
 AOI221_X1 _16368_ (.A(_07116_),
    .B1(_07117_),
    .B2(_06903_),
    .C1(_07062_),
    .C2(_07118_),
    .ZN(_07119_));
 AND2_X1 _16369_ (.A1(_14686_),
    .A2(_06233_),
    .ZN(_07120_));
 MUX2_X1 _16370_ (.A(net51),
    .B(_06907_),
    .S(_06931_),
    .Z(_07121_));
 AOI211_X2 _16371_ (.A(_06291_),
    .B(_07120_),
    .C1(_07121_),
    .C2(_06919_),
    .ZN(_07122_));
 AOI21_X4 _16372_ (.A(_14681_),
    .B1(_06965_),
    .B2(_06322_),
    .ZN(_07123_));
 MUX2_X1 _16373_ (.A(_06950_),
    .B(_07123_),
    .S(_06883_),
    .Z(_07124_));
 AOI21_X1 _16374_ (.A(_07122_),
    .B1(_07124_),
    .B2(_06293_),
    .ZN(_07125_));
 MUX2_X1 _16375_ (.A(_07119_),
    .B(_07125_),
    .S(_06278_),
    .Z(_07126_));
 MUX2_X1 _16376_ (.A(_07115_),
    .B(_07126_),
    .S(_00394_),
    .Z(_07127_));
 MUX2_X1 _16377_ (.A(_07100_),
    .B(_07127_),
    .S(_00393_),
    .Z(_00002_));
 MUX2_X1 _16378_ (.A(net64),
    .B(_06932_),
    .S(_06965_),
    .Z(_07128_));
 NAND2_X1 _16379_ (.A1(_06952_),
    .A2(_07128_),
    .ZN(_07129_));
 NAND2_X1 _16380_ (.A1(net64),
    .A2(_06917_),
    .ZN(_07130_));
 NAND3_X1 _16381_ (.A1(_07018_),
    .A2(_07041_),
    .A3(_07130_),
    .ZN(_07131_));
 AOI21_X1 _16382_ (.A(_06293_),
    .B1(_07129_),
    .B2(_07131_),
    .ZN(_07132_));
 NAND2_X1 _16383_ (.A1(_06953_),
    .A2(_07123_),
    .ZN(_07133_));
 OAI21_X1 _16384_ (.A(_07133_),
    .B1(_07022_),
    .B2(_06998_),
    .ZN(_07134_));
 AOI211_X2 _16385_ (.A(_00392_),
    .B(_07132_),
    .C1(_07134_),
    .C2(_06996_),
    .ZN(_07135_));
 NAND2_X1 _16386_ (.A1(net64),
    .A2(_06289_),
    .ZN(_07136_));
 NAND3_X1 _16387_ (.A1(_06965_),
    .A2(_06291_),
    .A3(_06870_),
    .ZN(_07137_));
 AOI21_X1 _16388_ (.A(_06919_),
    .B1(_07136_),
    .B2(_07137_),
    .ZN(_07138_));
 NAND2_X1 _16389_ (.A1(_06910_),
    .A2(_06289_),
    .ZN(_07139_));
 OAI21_X1 _16390_ (.A(_07139_),
    .B1(_07048_),
    .B2(_06903_),
    .ZN(_07140_));
 NAND2_X1 _16391_ (.A1(_07004_),
    .A2(_07062_),
    .ZN(_07141_));
 AOI221_X2 _16392_ (.A(_07138_),
    .B1(_07140_),
    .B2(_06883_),
    .C1(_07141_),
    .C2(_06323_),
    .ZN(_07142_));
 NAND3_X1 _16393_ (.A1(_06924_),
    .A2(_06238_),
    .A3(_07112_),
    .ZN(_07143_));
 AOI22_X1 _16394_ (.A1(_06890_),
    .A2(_06995_),
    .B1(_07112_),
    .B2(_06998_),
    .ZN(_07144_));
 OAI21_X1 _16395_ (.A(_07143_),
    .B1(_07144_),
    .B2(_06949_),
    .ZN(_07145_));
 NAND2_X2 _16396_ (.A1(net801),
    .A2(_06870_),
    .ZN(_07146_));
 AOI211_X2 _16397_ (.A(_06985_),
    .B(_07142_),
    .C1(_07145_),
    .C2(_07146_),
    .ZN(_07147_));
 NOR3_X1 _16398_ (.A1(_06929_),
    .A2(_07135_),
    .A3(_07147_),
    .ZN(_07148_));
 NOR2_X2 _16399_ (.A1(_06903_),
    .A2(_06917_),
    .ZN(_07149_));
 NAND3_X1 _16400_ (.A1(net43),
    .A2(_06952_),
    .A3(_06278_),
    .ZN(_07150_));
 INV_X2 _16401_ (.A(net1195),
    .ZN(_07151_));
 OAI21_X1 _16402_ (.A(_07150_),
    .B1(_06897_),
    .B2(_07151_),
    .ZN(_07152_));
 NOR2_X1 _16403_ (.A1(_06985_),
    .A2(_06293_),
    .ZN(_07153_));
 OAI22_X2 _16404_ (.A1(_06238_),
    .A2(_06954_),
    .B1(_07003_),
    .B2(_06935_),
    .ZN(_07154_));
 AOI221_X2 _16405_ (.A(_06596_),
    .B1(_07149_),
    .B2(_07152_),
    .C1(_07153_),
    .C2(_07154_),
    .ZN(_07155_));
 AOI21_X1 _16406_ (.A(_00390_),
    .B1(_07032_),
    .B2(_06956_),
    .ZN(_07156_));
 OAI21_X1 _16407_ (.A(_00391_),
    .B1(_07022_),
    .B2(_06998_),
    .ZN(_07157_));
 OAI21_X1 _16408_ (.A(_06985_),
    .B1(_07156_),
    .B2(_07157_),
    .ZN(_07158_));
 NAND2_X1 _16409_ (.A1(_06898_),
    .A2(_07024_),
    .ZN(_07159_));
 NAND3_X1 _16410_ (.A1(_00390_),
    .A2(_06925_),
    .A3(_06954_),
    .ZN(_07160_));
 AND3_X1 _16411_ (.A1(_06905_),
    .A2(_07159_),
    .A3(_07160_),
    .ZN(_07161_));
 OAI21_X1 _16412_ (.A(_07155_),
    .B1(_07158_),
    .B2(_07161_),
    .ZN(_07162_));
 NAND2_X1 _16413_ (.A1(_06874_),
    .A2(_07162_),
    .ZN(_07163_));
 MUX2_X1 _16414_ (.A(_06935_),
    .B(_06252_),
    .S(_06931_),
    .Z(_07164_));
 NAND2_X1 _16415_ (.A1(_07065_),
    .A2(_06925_),
    .ZN(_07165_));
 MUX2_X1 _16416_ (.A(_07016_),
    .B(_07165_),
    .S(_06291_),
    .Z(_07166_));
 AOI221_X2 _16417_ (.A(_06278_),
    .B1(_06887_),
    .B2(_07164_),
    .C1(_07166_),
    .C2(_06897_),
    .ZN(_07167_));
 OAI221_X1 _16418_ (.A(_07146_),
    .B1(_07021_),
    .B2(_07018_),
    .C1(_06961_),
    .C2(_07004_),
    .ZN(_07168_));
 MUX2_X2 _16419_ (.A(_06934_),
    .B(_06253_),
    .S(_06869_),
    .Z(_07169_));
 NOR2_X1 _16420_ (.A1(_06897_),
    .A2(_07169_),
    .ZN(_07170_));
 AOI21_X1 _16421_ (.A(_06948_),
    .B1(_06877_),
    .B2(_06925_),
    .ZN(_07171_));
 NOR2_X1 _16422_ (.A1(_07170_),
    .A2(_07171_),
    .ZN(_07172_));
 MUX2_X1 _16423_ (.A(_07168_),
    .B(_07172_),
    .S(_06293_),
    .Z(_07173_));
 AOI211_X2 _16424_ (.A(_00394_),
    .B(_07167_),
    .C1(_07173_),
    .C2(_00392_),
    .ZN(_07174_));
 NAND3_X1 _16425_ (.A1(_06925_),
    .A2(_07062_),
    .A3(_07032_),
    .ZN(_07175_));
 NAND2_X1 _16426_ (.A1(_06277_),
    .A2(_06596_),
    .ZN(_07176_));
 NOR2_X1 _16427_ (.A1(_06896_),
    .A2(_06932_),
    .ZN(_07177_));
 AOI21_X1 _16428_ (.A(_06292_),
    .B1(_07177_),
    .B2(_06915_),
    .ZN(_07178_));
 OAI21_X1 _16429_ (.A(_06877_),
    .B1(_14683_),
    .B2(_06935_),
    .ZN(_07179_));
 AOI221_X2 _16430_ (.A(_07176_),
    .B1(_07129_),
    .B2(_07178_),
    .C1(_07179_),
    .C2(_06942_),
    .ZN(_07180_));
 OAI221_X1 _16431_ (.A(_06982_),
    .B1(_06232_),
    .B2(_06219_),
    .C1(_06879_),
    .C2(_14678_),
    .ZN(_07181_));
 MUX2_X1 _16432_ (.A(_06915_),
    .B(_06890_),
    .S(_14683_),
    .Z(_07182_));
 NAND2_X1 _16433_ (.A1(_00390_),
    .A2(_07182_),
    .ZN(_07183_));
 NAND3_X1 _16434_ (.A1(_06905_),
    .A2(_07181_),
    .A3(_07183_),
    .ZN(_07184_));
 NAND2_X1 _16435_ (.A1(_06278_),
    .A2(_06596_),
    .ZN(_07185_));
 NOR2_X1 _16436_ (.A1(_06899_),
    .A2(_06900_),
    .ZN(_07186_));
 AOI221_X1 _16437_ (.A(_07185_),
    .B1(_07062_),
    .B2(_07186_),
    .C1(_06944_),
    .C2(_07041_),
    .ZN(_07187_));
 AOI22_X1 _16438_ (.A1(_07175_),
    .A2(_07180_),
    .B1(_07184_),
    .B2(_07187_),
    .ZN(_07188_));
 NAND2_X1 _16439_ (.A1(_00393_),
    .A2(_07188_),
    .ZN(_07189_));
 OAI22_X1 _16440_ (.A1(_07148_),
    .A2(_07163_),
    .B1(_07174_),
    .B2(_07189_),
    .ZN(_00003_));
 MUX2_X1 _16441_ (.A(_06253_),
    .B(_06880_),
    .S(_14669_),
    .Z(_07190_));
 MUX2_X1 _16442_ (.A(_07164_),
    .B(_07190_),
    .S(_06896_),
    .Z(_07191_));
 OAI21_X1 _16443_ (.A(_06895_),
    .B1(_06960_),
    .B2(_06948_),
    .ZN(_07192_));
 MUX2_X1 _16444_ (.A(_07191_),
    .B(_07192_),
    .S(_06904_),
    .Z(_07193_));
 MUX2_X2 _16445_ (.A(_06934_),
    .B(_06868_),
    .S(_06931_),
    .Z(_07194_));
 MUX2_X1 _16446_ (.A(_06982_),
    .B(_07194_),
    .S(_06292_),
    .Z(_07195_));
 NAND2_X1 _16447_ (.A1(_06949_),
    .A2(_07195_),
    .ZN(_07196_));
 NAND3_X1 _16448_ (.A1(net65),
    .A2(_06292_),
    .A3(_06323_),
    .ZN(_07197_));
 OAI21_X1 _16449_ (.A(_07197_),
    .B1(_06995_),
    .B2(_06879_),
    .ZN(_07198_));
 AOI21_X1 _16450_ (.A(_06985_),
    .B1(_07198_),
    .B2(_06953_),
    .ZN(_07199_));
 AOI22_X1 _16451_ (.A1(_06985_),
    .A2(_07193_),
    .B1(_07196_),
    .B2(_07199_),
    .ZN(_07200_));
 NOR2_X1 _16452_ (.A1(_06289_),
    .A2(_06322_),
    .ZN(_07201_));
 AOI22_X2 _16453_ (.A1(_07035_),
    .A2(_06884_),
    .B1(_07201_),
    .B2(_06970_),
    .ZN(_07202_));
 AOI22_X1 _16454_ (.A1(net65),
    .A2(_07112_),
    .B1(_07201_),
    .B2(_06998_),
    .ZN(_07203_));
 NOR2_X2 _16455_ (.A1(_06291_),
    .A2(_06322_),
    .ZN(_07204_));
 AOI21_X1 _16456_ (.A(_07149_),
    .B1(_07204_),
    .B2(_06948_),
    .ZN(_07205_));
 OAI221_X1 _16457_ (.A(_07202_),
    .B1(_07203_),
    .B2(_06897_),
    .C1(_06935_),
    .C2(_07205_),
    .ZN(_07206_));
 MUX2_X1 _16458_ (.A(_06959_),
    .B(net42),
    .S(net999),
    .Z(_07207_));
 MUX2_X1 _16459_ (.A(_07090_),
    .B(_07207_),
    .S(_06236_),
    .Z(_07208_));
 MUX2_X1 _16460_ (.A(_06907_),
    .B(net42),
    .S(_06916_),
    .Z(_07209_));
 MUX2_X1 _16461_ (.A(_07088_),
    .B(_07209_),
    .S(_06919_),
    .Z(_07210_));
 MUX2_X1 _16462_ (.A(_07208_),
    .B(_07210_),
    .S(_06292_),
    .Z(_07211_));
 MUX2_X1 _16463_ (.A(_07206_),
    .B(_07211_),
    .S(_06985_),
    .Z(_07212_));
 MUX2_X1 _16464_ (.A(_07200_),
    .B(_07212_),
    .S(_00394_),
    .Z(_07213_));
 MUX2_X1 _16465_ (.A(_07004_),
    .B(net66),
    .S(_06881_),
    .Z(_07214_));
 AOI22_X1 _16466_ (.A1(_06924_),
    .A2(_07204_),
    .B1(_07214_),
    .B2(_06995_),
    .ZN(_07215_));
 NOR2_X1 _16467_ (.A1(_06949_),
    .A2(_07215_),
    .ZN(_07216_));
 AOI21_X1 _16468_ (.A(_06596_),
    .B1(_07112_),
    .B2(net801),
    .ZN(_07217_));
 AOI21_X1 _16469_ (.A(_07112_),
    .B1(_07012_),
    .B2(_06995_),
    .ZN(_07218_));
 OAI21_X1 _16470_ (.A(_07217_),
    .B1(_07218_),
    .B2(_06898_),
    .ZN(_07219_));
 AOI21_X1 _16471_ (.A(_07149_),
    .B1(_06887_),
    .B2(net1000),
    .ZN(_07220_));
 OAI21_X1 _16472_ (.A(_00394_),
    .B1(_07220_),
    .B2(net66),
    .ZN(_07221_));
 AOI221_X1 _16473_ (.A(_06896_),
    .B1(net64),
    .B2(_07112_),
    .C1(_07201_),
    .C2(_07004_),
    .ZN(_07222_));
 AOI22_X1 _16474_ (.A1(_14659_),
    .A2(_06989_),
    .B1(_07204_),
    .B2(net66),
    .ZN(_07223_));
 AOI21_X1 _16475_ (.A(_07222_),
    .B1(_07223_),
    .B2(_06953_),
    .ZN(_07224_));
 OAI22_X1 _16476_ (.A1(_07216_),
    .A2(_07219_),
    .B1(_07221_),
    .B2(_07224_),
    .ZN(_07225_));
 NAND2_X1 _16477_ (.A1(_06910_),
    .A2(_06323_),
    .ZN(_07226_));
 AOI21_X1 _16478_ (.A(_06948_),
    .B1(_07048_),
    .B2(_07226_),
    .ZN(_07227_));
 MUX2_X1 _16479_ (.A(net1195),
    .B(_06971_),
    .S(_06237_),
    .Z(_07228_));
 NAND2_X1 _16480_ (.A1(_06293_),
    .A2(_14678_),
    .ZN(_07229_));
 OAI221_X1 _16481_ (.A(_06929_),
    .B1(_06988_),
    .B2(_07227_),
    .C1(_07228_),
    .C2(_07229_),
    .ZN(_07230_));
 NOR2_X1 _16482_ (.A1(_06934_),
    .A2(_06323_),
    .ZN(_07231_));
 OAI221_X1 _16483_ (.A(_06995_),
    .B1(_14678_),
    .B2(_07151_),
    .C1(_07231_),
    .C2(_06897_),
    .ZN(_07232_));
 NAND2_X1 _16484_ (.A1(_06886_),
    .A2(_06917_),
    .ZN(_07233_));
 INV_X1 _16485_ (.A(_14690_),
    .ZN(_07234_));
 OAI221_X1 _16486_ (.A(_06954_),
    .B1(_07233_),
    .B2(_07004_),
    .C1(_06953_),
    .C2(_07234_),
    .ZN(_07235_));
 OAI21_X1 _16487_ (.A(_07232_),
    .B1(_07235_),
    .B2(_06996_),
    .ZN(_07236_));
 OAI21_X1 _16488_ (.A(_07230_),
    .B1(_07236_),
    .B2(_06929_),
    .ZN(_07237_));
 MUX2_X1 _16489_ (.A(_07225_),
    .B(_07237_),
    .S(_00392_),
    .Z(_07238_));
 MUX2_X1 _16490_ (.A(_07213_),
    .B(_07238_),
    .S(_00393_),
    .Z(_00004_));
 NAND3_X1 _16491_ (.A1(net801),
    .A2(net66),
    .A3(_06293_),
    .ZN(_07239_));
 NAND2_X1 _16492_ (.A1(_06903_),
    .A2(_06881_),
    .ZN(_07240_));
 OAI21_X1 _16493_ (.A(_07239_),
    .B1(_07240_),
    .B2(net66),
    .ZN(_07241_));
 OAI21_X1 _16494_ (.A(_07136_),
    .B1(_07016_),
    .B2(_06904_),
    .ZN(_07242_));
 MUX2_X1 _16495_ (.A(_07241_),
    .B(_07242_),
    .S(_00390_),
    .Z(_07243_));
 AOI21_X1 _16496_ (.A(net801),
    .B1(_07233_),
    .B2(_07136_),
    .ZN(_07244_));
 OR2_X1 _16497_ (.A1(_00393_),
    .A2(_07244_),
    .ZN(_07245_));
 AOI21_X1 _16498_ (.A(_06996_),
    .B1(_06940_),
    .B2(_06989_),
    .ZN(_07246_));
 AND3_X1 _16499_ (.A1(_06996_),
    .A2(_06933_),
    .A3(_06936_),
    .ZN(_07247_));
 OAI21_X1 _16500_ (.A(_06898_),
    .B1(_07246_),
    .B2(_07247_),
    .ZN(_07248_));
 NOR3_X1 _16501_ (.A1(_06969_),
    .A2(_07149_),
    .A3(_07204_),
    .ZN(_07249_));
 AOI221_X2 _16502_ (.A(_07249_),
    .B1(_07149_),
    .B2(net1000),
    .C1(_14662_),
    .C2(_07204_),
    .ZN(_07250_));
 OAI21_X1 _16503_ (.A(_07248_),
    .B1(_07250_),
    .B2(_06898_),
    .ZN(_07251_));
 OAI221_X1 _16504_ (.A(_06930_),
    .B1(_07243_),
    .B2(_07245_),
    .C1(_07251_),
    .C2(_06874_),
    .ZN(_07252_));
 NAND2_X1 _16505_ (.A1(net1000),
    .A2(_06584_),
    .ZN(_07253_));
 OAI21_X1 _16506_ (.A(_07253_),
    .B1(_06584_),
    .B2(_06879_),
    .ZN(_07254_));
 OAI221_X2 _16507_ (.A(_06953_),
    .B1(_06585_),
    .B2(_06918_),
    .C1(_07254_),
    .C2(_14678_),
    .ZN(_07255_));
 NAND2_X1 _16508_ (.A1(_06873_),
    .A2(_06900_),
    .ZN(_07256_));
 NAND3_X1 _16509_ (.A1(_06238_),
    .A2(_07253_),
    .A3(_07256_),
    .ZN(_07257_));
 AOI221_X2 _16510_ (.A(_06996_),
    .B1(_06585_),
    .B2(_06899_),
    .C1(_07255_),
    .C2(_07257_),
    .ZN(_07258_));
 AOI21_X1 _16511_ (.A(_07033_),
    .B1(_07177_),
    .B2(_06924_),
    .ZN(_07259_));
 MUX2_X1 _16512_ (.A(_06978_),
    .B(net65),
    .S(_06870_),
    .Z(_07260_));
 MUX2_X1 _16513_ (.A(_07194_),
    .B(_07260_),
    .S(_06238_),
    .Z(_07261_));
 MUX2_X1 _16514_ (.A(_07259_),
    .B(_07261_),
    .S(_00393_),
    .Z(_07262_));
 AOI21_X1 _16515_ (.A(_07258_),
    .B1(_07262_),
    .B2(_00391_),
    .ZN(_07263_));
 NAND2_X1 _16516_ (.A1(_06278_),
    .A2(_06595_),
    .ZN(_07264_));
 MUX2_X1 _16517_ (.A(_06978_),
    .B(_06924_),
    .S(_06916_),
    .Z(_07265_));
 MUX2_X1 _16518_ (.A(_06876_),
    .B(_06890_),
    .S(_06880_),
    .Z(_07266_));
 MUX2_X1 _16519_ (.A(_07265_),
    .B(_07266_),
    .S(_06919_),
    .Z(_07267_));
 AOI21_X1 _16520_ (.A(_06919_),
    .B1(_06932_),
    .B2(_06879_),
    .ZN(_07268_));
 AOI21_X1 _16521_ (.A(_07268_),
    .B1(_06948_),
    .B2(_06955_),
    .ZN(_07269_));
 MUX2_X1 _16522_ (.A(_07267_),
    .B(_07269_),
    .S(_06986_),
    .Z(_07270_));
 MUX2_X1 _16523_ (.A(_06924_),
    .B(_06879_),
    .S(_06932_),
    .Z(_07271_));
 OAI221_X1 _16524_ (.A(_06995_),
    .B1(_07022_),
    .B2(_06890_),
    .C1(_07271_),
    .C2(_07018_),
    .ZN(_07272_));
 NOR2_X1 _16525_ (.A1(_06920_),
    .A2(_07028_),
    .ZN(_07273_));
 OAI21_X1 _16526_ (.A(_07272_),
    .B1(_07273_),
    .B2(_06988_),
    .ZN(_07274_));
 MUX2_X1 _16527_ (.A(_07270_),
    .B(_07274_),
    .S(_06585_),
    .Z(_07275_));
 OAI221_X1 _16528_ (.A(_06585_),
    .B1(_06911_),
    .B2(_06948_),
    .C1(_14683_),
    .C2(_06915_),
    .ZN(_07276_));
 MUX2_X1 _16529_ (.A(_07151_),
    .B(net66),
    .S(_06932_),
    .Z(_07277_));
 OAI221_X1 _16530_ (.A(_06873_),
    .B1(_07022_),
    .B2(net43),
    .C1(_07277_),
    .C2(_07018_),
    .ZN(_07278_));
 AND3_X1 _16531_ (.A1(_06996_),
    .A2(_07276_),
    .A3(_07278_),
    .ZN(_07279_));
 MUX2_X1 _16532_ (.A(net43),
    .B(_06959_),
    .S(_06870_),
    .Z(_07280_));
 AOI221_X2 _16533_ (.A(_06584_),
    .B1(_07002_),
    .B2(_14662_),
    .C1(_07280_),
    .C2(_06237_),
    .ZN(_07281_));
 OAI22_X1 _16534_ (.A1(_06998_),
    .A2(_07070_),
    .B1(_07169_),
    .B2(_06953_),
    .ZN(_07282_));
 AOI21_X1 _16535_ (.A(_07281_),
    .B1(_07282_),
    .B2(_00393_),
    .ZN(_07283_));
 AOI21_X1 _16536_ (.A(_07279_),
    .B1(_07283_),
    .B2(_06905_),
    .ZN(_07284_));
 MUX2_X1 _16537_ (.A(_07275_),
    .B(_07284_),
    .S(_00394_),
    .Z(_07285_));
 OAI221_X2 _16538_ (.A(_07252_),
    .B1(_07263_),
    .B2(_07264_),
    .C1(_07285_),
    .C2(_00392_),
    .ZN(_00005_));
 MUX2_X1 _16539_ (.A(_07090_),
    .B(_07194_),
    .S(_06292_),
    .Z(_07286_));
 OAI221_X2 _16540_ (.A(_06873_),
    .B1(_06938_),
    .B2(_06943_),
    .C1(_07286_),
    .C2(_06898_),
    .ZN(_07287_));
 AND2_X1 _16541_ (.A1(_07018_),
    .A2(_07169_),
    .ZN(_07288_));
 OAI21_X1 _16542_ (.A(_06904_),
    .B1(_07070_),
    .B2(net43),
    .ZN(_07289_));
 OAI21_X1 _16543_ (.A(_06585_),
    .B1(_07288_),
    .B2(_07289_),
    .ZN(_07290_));
 INV_X1 _16544_ (.A(_14679_),
    .ZN(_07291_));
 AOI221_X2 _16545_ (.A(_06986_),
    .B1(_06918_),
    .B2(_06921_),
    .C1(_06948_),
    .C2(_07291_),
    .ZN(_07292_));
 OAI21_X1 _16546_ (.A(_07287_),
    .B1(_07290_),
    .B2(_07292_),
    .ZN(_07293_));
 MUX2_X1 _16547_ (.A(_14662_),
    .B(_06934_),
    .S(_06319_),
    .Z(_07294_));
 MUX2_X1 _16548_ (.A(_14676_),
    .B(_06971_),
    .S(_06869_),
    .Z(_07295_));
 MUX2_X1 _16549_ (.A(_07294_),
    .B(_07295_),
    .S(_06236_),
    .Z(_07296_));
 MUX2_X1 _16550_ (.A(_06907_),
    .B(_06253_),
    .S(_06869_),
    .Z(_07297_));
 MUX2_X1 _16551_ (.A(_06876_),
    .B(_06253_),
    .S(_06321_),
    .Z(_07298_));
 MUX2_X1 _16552_ (.A(_07297_),
    .B(_07298_),
    .S(_06886_),
    .Z(_07299_));
 MUX2_X1 _16553_ (.A(_07296_),
    .B(_07299_),
    .S(_06873_),
    .Z(_07300_));
 MUX2_X1 _16554_ (.A(_07169_),
    .B(_07298_),
    .S(_06886_),
    .Z(_07301_));
 MUX2_X1 _16555_ (.A(net1193),
    .B(_06265_),
    .S(_06916_),
    .Z(_07302_));
 OAI22_X1 _16556_ (.A1(_06890_),
    .A2(_07233_),
    .B1(_07302_),
    .B2(_06896_),
    .ZN(_07303_));
 MUX2_X1 _16557_ (.A(_07301_),
    .B(_07303_),
    .S(_06873_),
    .Z(_07304_));
 MUX2_X1 _16558_ (.A(_07300_),
    .B(_07304_),
    .S(_06293_),
    .Z(_07305_));
 MUX2_X1 _16559_ (.A(_07293_),
    .B(_07305_),
    .S(_00394_),
    .Z(_07306_));
 NOR2_X1 _16560_ (.A1(_14662_),
    .A2(_07070_),
    .ZN(_07307_));
 OAI21_X1 _16561_ (.A(_07146_),
    .B1(_06894_),
    .B2(_06953_),
    .ZN(_07308_));
 NOR3_X1 _16562_ (.A1(_06873_),
    .A2(_07307_),
    .A3(_07308_),
    .ZN(_07309_));
 AOI21_X1 _16563_ (.A(_06237_),
    .B1(net801),
    .B2(_06870_),
    .ZN(_07310_));
 AOI211_X2 _16564_ (.A(_06585_),
    .B(_07310_),
    .C1(_07265_),
    .C2(_06238_),
    .ZN(_07311_));
 NOR3_X1 _16565_ (.A1(_06905_),
    .A2(_07309_),
    .A3(_07311_),
    .ZN(_07312_));
 NOR2_X1 _16566_ (.A1(_14680_),
    .A2(_06952_),
    .ZN(_07313_));
 AOI21_X1 _16567_ (.A(_07313_),
    .B1(_07194_),
    .B2(_06953_),
    .ZN(_07314_));
 AND2_X1 _16568_ (.A1(_06949_),
    .A2(_07128_),
    .ZN(_07315_));
 OAI221_X1 _16569_ (.A(_06585_),
    .B1(_06918_),
    .B2(_06238_),
    .C1(_14669_),
    .C2(_14678_),
    .ZN(_07316_));
 OAI221_X1 _16570_ (.A(_06905_),
    .B1(_00393_),
    .B2(_07314_),
    .C1(_07315_),
    .C2(_07316_),
    .ZN(_07317_));
 NAND2_X1 _16571_ (.A1(_06929_),
    .A2(_07317_),
    .ZN(_07318_));
 NAND2_X1 _16572_ (.A1(_06919_),
    .A2(_14659_),
    .ZN(_07319_));
 AOI221_X1 _16573_ (.A(_06583_),
    .B1(_06997_),
    .B2(_06919_),
    .C1(_07319_),
    .C2(net66),
    .ZN(_07320_));
 MUX2_X1 _16574_ (.A(_06876_),
    .B(net1195),
    .S(_06917_),
    .Z(_07321_));
 MUX2_X1 _16575_ (.A(_06991_),
    .B(_07321_),
    .S(_06952_),
    .Z(_07322_));
 AOI21_X1 _16576_ (.A(_07320_),
    .B1(_07322_),
    .B2(_06873_),
    .ZN(_07323_));
 NAND2_X1 _16577_ (.A1(net1195),
    .A2(_06870_),
    .ZN(_07324_));
 AOI21_X1 _16578_ (.A(_06897_),
    .B1(_07102_),
    .B2(_07324_),
    .ZN(_07325_));
 OR2_X1 _16579_ (.A1(_06873_),
    .A2(_07084_),
    .ZN(_07326_));
 INV_X1 _16580_ (.A(_14684_),
    .ZN(_07327_));
 MUX2_X1 _16581_ (.A(_07327_),
    .B(_07260_),
    .S(_06952_),
    .Z(_07328_));
 OAI22_X1 _16582_ (.A1(_07325_),
    .A2(_07326_),
    .B1(_07328_),
    .B2(_06585_),
    .ZN(_07329_));
 MUX2_X1 _16583_ (.A(_07323_),
    .B(_07329_),
    .S(_06996_),
    .Z(_07330_));
 OAI22_X1 _16584_ (.A1(_07312_),
    .A2(_07318_),
    .B1(_07330_),
    .B2(_06929_),
    .ZN(_07331_));
 MUX2_X1 _16585_ (.A(_07306_),
    .B(_07331_),
    .S(_00392_),
    .Z(_00006_));
 NOR2_X1 _16586_ (.A1(_07151_),
    .A2(_07018_),
    .ZN(_07332_));
 OAI21_X1 _16587_ (.A(_06870_),
    .B1(net1205),
    .B2(_06952_),
    .ZN(_07333_));
 OAI221_X2 _16588_ (.A(_06904_),
    .B1(_07332_),
    .B2(_07333_),
    .C1(_14678_),
    .C2(_06959_),
    .ZN(_07334_));
 NOR2_X1 _16589_ (.A1(_06897_),
    .A2(_07190_),
    .ZN(_07335_));
 OAI21_X1 _16590_ (.A(_06996_),
    .B1(_06970_),
    .B2(_07335_),
    .ZN(_07336_));
 AOI21_X1 _16591_ (.A(_07176_),
    .B1(_07334_),
    .B2(_07336_),
    .ZN(_07337_));
 NOR3_X1 _16592_ (.A1(_06235_),
    .A2(_06291_),
    .A3(_07294_),
    .ZN(_07338_));
 OR3_X1 _16593_ (.A1(_06278_),
    .A2(_06596_),
    .A3(_07338_),
    .ZN(_07339_));
 INV_X1 _16594_ (.A(_07003_),
    .ZN(_07340_));
 OAI222_X2 _16595_ (.A1(_06237_),
    .A2(_06913_),
    .B1(_06961_),
    .B2(_14662_),
    .C1(net51),
    .C2(_07340_),
    .ZN(_07341_));
 AOI221_X2 _16596_ (.A(_07339_),
    .B1(_07123_),
    .B2(_06887_),
    .C1(_06995_),
    .C2(_07341_),
    .ZN(_07342_));
 AOI21_X1 _16597_ (.A(_06938_),
    .B1(_06933_),
    .B2(_06913_),
    .ZN(_07343_));
 NAND2_X1 _16598_ (.A1(_06882_),
    .A2(_07049_),
    .ZN(_07344_));
 AOI21_X1 _16599_ (.A(_07343_),
    .B1(_07344_),
    .B2(_07062_),
    .ZN(_07345_));
 NOR2_X1 _16600_ (.A1(_06952_),
    .A2(_07194_),
    .ZN(_07346_));
 OAI21_X1 _16601_ (.A(_06986_),
    .B1(_07307_),
    .B2(_07346_),
    .ZN(_07347_));
 AND3_X1 _16602_ (.A1(_06872_),
    .A2(_07345_),
    .A3(_07347_),
    .ZN(_07348_));
 MUX2_X1 _16603_ (.A(_07004_),
    .B(_06868_),
    .S(_06291_),
    .Z(_07349_));
 AOI22_X1 _16604_ (.A1(_06879_),
    .A2(_07204_),
    .B1(_07349_),
    .B2(_06323_),
    .ZN(_07350_));
 NOR2_X1 _16605_ (.A1(_07018_),
    .A2(_07350_),
    .ZN(_07351_));
 NAND2_X1 _16606_ (.A1(_06237_),
    .A2(_06986_),
    .ZN(_07352_));
 AOI21_X1 _16607_ (.A(_07352_),
    .B1(_06943_),
    .B2(_07041_),
    .ZN(_07353_));
 AOI22_X1 _16608_ (.A1(_06879_),
    .A2(_07002_),
    .B1(_07164_),
    .B2(_06883_),
    .ZN(_07354_));
 NOR2_X1 _16609_ (.A1(_06986_),
    .A2(_07354_),
    .ZN(_07355_));
 NOR4_X1 _16610_ (.A1(_07185_),
    .A2(_07351_),
    .A3(_07353_),
    .A4(_07355_),
    .ZN(_07356_));
 OR4_X1 _16611_ (.A1(_07337_),
    .A2(_07342_),
    .A3(_07348_),
    .A4(_07356_),
    .ZN(_07357_));
 OAI221_X2 _16612_ (.A(_06897_),
    .B1(_06986_),
    .B2(_07302_),
    .C1(_07240_),
    .C2(_07151_),
    .ZN(_07358_));
 NAND2_X1 _16613_ (.A1(_06292_),
    .A2(_06989_),
    .ZN(_07359_));
 OAI221_X1 _16614_ (.A(_07018_),
    .B1(_06911_),
    .B2(_07359_),
    .C1(_06995_),
    .C2(_06879_),
    .ZN(_07360_));
 AOI21_X1 _16615_ (.A(_07185_),
    .B1(_07358_),
    .B2(_07360_),
    .ZN(_07361_));
 NAND3_X1 _16616_ (.A1(_06882_),
    .A2(_06884_),
    .A3(_07032_),
    .ZN(_07362_));
 MUX2_X1 _16617_ (.A(_06965_),
    .B(_06920_),
    .S(_06235_),
    .Z(_07363_));
 OAI21_X1 _16618_ (.A(_07130_),
    .B1(_07067_),
    .B2(_06291_),
    .ZN(_07364_));
 AOI221_X1 _16619_ (.A(_07264_),
    .B1(_07363_),
    .B2(_06292_),
    .C1(_07364_),
    .C2(_06237_),
    .ZN(_07365_));
 AOI21_X1 _16620_ (.A(_14686_),
    .B1(_06252_),
    .B2(_06916_),
    .ZN(_07366_));
 MUX2_X1 _16621_ (.A(_07105_),
    .B(_07366_),
    .S(_06886_),
    .Z(_07367_));
 MUX2_X1 _16622_ (.A(_14661_),
    .B(_06935_),
    .S(_06321_),
    .Z(_07368_));
 MUX2_X1 _16623_ (.A(_07234_),
    .B(_07368_),
    .S(_06886_),
    .Z(_07369_));
 MUX2_X1 _16624_ (.A(_07367_),
    .B(_07369_),
    .S(_06903_),
    .Z(_07370_));
 NOR2_X1 _16625_ (.A1(_06887_),
    .A2(_07002_),
    .ZN(_07371_));
 AOI22_X1 _16626_ (.A1(_06998_),
    .A2(_06896_),
    .B1(_07062_),
    .B2(_06915_),
    .ZN(_07372_));
 OAI221_X1 _16627_ (.A(_07240_),
    .B1(_07371_),
    .B2(_06971_),
    .C1(_07372_),
    .C2(_06870_),
    .ZN(_07373_));
 MUX2_X1 _16628_ (.A(_07370_),
    .B(_07373_),
    .S(_06929_),
    .Z(_07374_));
 AOI221_X2 _16629_ (.A(_07361_),
    .B1(_07362_),
    .B2(_07365_),
    .C1(_06985_),
    .C2(_07374_),
    .ZN(_07375_));
 MUX2_X1 _16630_ (.A(_07357_),
    .B(_07375_),
    .S(_06874_),
    .Z(_00007_));
 BUF_X8 _16631_ (.A(_06475_),
    .Z(_07376_));
 BUF_X16 _16632_ (.A(_07376_),
    .Z(_07377_));
 BUF_X16 _16633_ (.A(_07377_),
    .Z(_14692_));
 BUF_X8 _16634_ (.A(_06503_),
    .Z(_07378_));
 BUF_X8 _16635_ (.A(_07378_),
    .Z(_07379_));
 BUF_X8 _16636_ (.A(_07379_),
    .Z(_07380_));
 BUF_X8 _16637_ (.A(_07380_),
    .Z(_14712_));
 BUF_X8 _16638_ (.A(_06461_),
    .Z(_07381_));
 BUF_X16 _16639_ (.A(_07381_),
    .Z(_14693_));
 BUF_X4 _16640_ (.A(_06550_),
    .Z(_07382_));
 BUF_X4 _16641_ (.A(_14708_),
    .Z(_07383_));
 CLKBUF_X3 _16642_ (.A(_06509_),
    .Z(_07384_));
 BUF_X4 _16643_ (.A(_06521_),
    .Z(_07385_));
 NAND3_X1 _16644_ (.A1(_07383_),
    .A2(_07384_),
    .A3(_07385_),
    .ZN(_07386_));
 CLKBUF_X3 _16645_ (.A(_14699_),
    .Z(_07387_));
 NOR2_X4 _16646_ (.A1(_06266_),
    .A2(net52),
    .ZN(_07388_));
 BUF_X4 _16647_ (.A(_07388_),
    .Z(_07389_));
 NOR2_X1 _16648_ (.A1(net18),
    .A2(_06514_),
    .ZN(_07390_));
 NOR2_X1 _16649_ (.A1(net18),
    .A2(_06512_),
    .ZN(_07391_));
 MUX2_X1 _16650_ (.A(_07390_),
    .B(_07391_),
    .S(_06519_),
    .Z(_07392_));
 BUF_X4 _16651_ (.A(_07392_),
    .Z(_07393_));
 BUF_X4 _16652_ (.A(_07393_),
    .Z(_07394_));
 OAI21_X2 _16653_ (.A(_07387_),
    .B1(_07389_),
    .B2(_07394_),
    .ZN(_07395_));
 NAND3_X2 _16654_ (.A1(_06506_),
    .A2(_07386_),
    .A3(_07395_),
    .ZN(_07396_));
 NOR4_X4 _16655_ (.A1(_06449_),
    .A2(net1236),
    .A3(_07388_),
    .A4(_07393_),
    .ZN(_07397_));
 OR2_X1 _16656_ (.A1(_06267_),
    .A2(net214),
    .ZN(_07398_));
 NAND2_X1 _16657_ (.A1(_06266_),
    .A2(_06454_),
    .ZN(_07399_));
 NAND2_X1 _16658_ (.A1(_06266_),
    .A2(_06452_),
    .ZN(_07400_));
 MUX2_X2 _16659_ (.A(_07399_),
    .B(_07400_),
    .S(_06459_),
    .Z(_07401_));
 AOI22_X4 _16660_ (.A1(_07398_),
    .A2(_07401_),
    .B1(_06509_),
    .B2(_06521_),
    .ZN(_07402_));
 OAI21_X1 _16661_ (.A(_07379_),
    .B1(_07397_),
    .B2(_07402_),
    .ZN(_07403_));
 AND3_X1 _16662_ (.A1(_07382_),
    .A2(_07396_),
    .A3(_07403_),
    .ZN(_07404_));
 NOR2_X4 _16663_ (.A1(_06504_),
    .A2(_06522_),
    .ZN(_07405_));
 CLKBUF_X1 hold776 (.A(net226),
    .Z(net1239));
 BUF_X4 _16665_ (.A(_14706_),
    .Z(_07407_));
 BUF_X8 clone66 (.A(_06868_),
    .Z(net66));
 OAI21_X2 _16667_ (.A(_14710_),
    .B1(_07388_),
    .B2(_07393_),
    .ZN(_07409_));
 BUF_X4 _16668_ (.A(_06522_),
    .Z(_07410_));
 OAI21_X1 _16669_ (.A(_07409_),
    .B1(_07410_),
    .B2(_07387_),
    .ZN(_07411_));
 BUF_X4 _16670_ (.A(_06505_),
    .Z(_07412_));
 AOI221_X1 _16671_ (.A(_06550_),
    .B1(_07405_),
    .B2(_07407_),
    .C1(_07411_),
    .C2(_07412_),
    .ZN(_07413_));
 NOR3_X1 _16672_ (.A1(_06540_),
    .A2(_07404_),
    .A3(_07413_),
    .ZN(_07414_));
 CLKBUF_X3 _16673_ (.A(_06537_),
    .Z(_07415_));
 CLKBUF_X3 _16674_ (.A(_07415_),
    .Z(_07416_));
 CLKBUF_X3 _16675_ (.A(_07416_),
    .Z(_07417_));
 NOR2_X1 _16676_ (.A1(_06504_),
    .A2(_06523_),
    .ZN(_07418_));
 BUF_X4 _16677_ (.A(_07418_),
    .Z(_07419_));
 BUF_X8 clone18 (.A(_06226_),
    .Z(net18));
 INV_X1 _16679_ (.A(_14704_),
    .ZN(_07421_));
 NAND3_X1 _16680_ (.A1(_14710_),
    .A2(_07384_),
    .A3(_07385_),
    .ZN(_07422_));
 BUF_X8 _16681_ (.A(_07387_),
    .Z(_07423_));
 OAI21_X1 _16682_ (.A(_07422_),
    .B1(_06524_),
    .B2(_07423_),
    .ZN(_07424_));
 AOI221_X1 _16683_ (.A(_06550_),
    .B1(_07419_),
    .B2(_07421_),
    .C1(_07424_),
    .C2(_07412_),
    .ZN(_07425_));
 BUF_X4 _16684_ (.A(_14695_),
    .Z(_07426_));
 BUF_X8 _16685_ (.A(_07426_),
    .Z(_07427_));
 BUF_X4 _16686_ (.A(_06524_),
    .Z(_07428_));
 AOI221_X1 _16687_ (.A(_06551_),
    .B1(_07419_),
    .B2(_07427_),
    .C1(_14720_),
    .C2(_07428_),
    .ZN(_07429_));
 NOR3_X1 _16688_ (.A1(_07417_),
    .A2(_07425_),
    .A3(_07429_),
    .ZN(_07430_));
 OR2_X1 _16689_ (.A1(_07414_),
    .A2(_07430_),
    .ZN(_07431_));
 NAND3_X4 _16690_ (.A1(_14704_),
    .A2(_06509_),
    .A3(_06521_),
    .ZN(_07432_));
 INV_X8 _16691_ (.A(_07426_),
    .ZN(_07433_));
 OAI21_X4 _16692_ (.A(_07433_),
    .B1(_07388_),
    .B2(_07393_),
    .ZN(_07434_));
 NAND3_X4 _16693_ (.A1(_06506_),
    .A2(_07432_),
    .A3(net1051),
    .ZN(_07435_));
 NOR2_X2 clone28 (.A1(_06350_),
    .A2(_06338_),
    .ZN(net28));
 OAI21_X2 _16695_ (.A(_14694_),
    .B1(_07389_),
    .B2(_07394_),
    .ZN(_07437_));
 NAND3_X1 _16696_ (.A1(_07379_),
    .A2(_07386_),
    .A3(_07437_),
    .ZN(_07438_));
 NAND2_X2 _16697_ (.A1(_07438_),
    .A2(_07435_),
    .ZN(_07439_));
 NOR3_X4 _16698_ (.A1(_07426_),
    .A2(_06503_),
    .A3(_06522_),
    .ZN(_07440_));
 XNOR2_X2 _16699_ (.A(_06503_),
    .B(_06523_),
    .ZN(_07441_));
 AOI221_X1 _16700_ (.A(_07440_),
    .B1(_07441_),
    .B2(net956),
    .C1(_14704_),
    .C2(_07418_),
    .ZN(_07442_));
 MUX2_X1 _16701_ (.A(_07439_),
    .B(_07442_),
    .S(_07382_),
    .Z(_07443_));
 CLKBUF_X3 _16702_ (.A(_07412_),
    .Z(_07444_));
 NOR2_X2 _16703_ (.A1(_06524_),
    .A2(_06551_),
    .ZN(_07445_));
 NAND3_X1 _16704_ (.A1(_07427_),
    .A2(_07444_),
    .A3(_07445_),
    .ZN(_07446_));
 CLKBUF_X3 _16705_ (.A(_07410_),
    .Z(_07447_));
 NOR3_X4 _16706_ (.A1(_07427_),
    .A2(_07388_),
    .A3(_07393_),
    .ZN(_07448_));
 AOI22_X2 _16707_ (.A1(_07377_),
    .A2(_07447_),
    .B1(_07448_),
    .B2(_07382_),
    .ZN(_07449_));
 XNOR2_X2 _16708_ (.A(net1225),
    .B(_06523_),
    .ZN(_07450_));
 MUX2_X1 _16709_ (.A(_07441_),
    .B(_07450_),
    .S(_06463_),
    .Z(_07451_));
 CLKBUF_X3 _16710_ (.A(_07382_),
    .Z(_07452_));
 OAI221_X1 _16711_ (.A(_07446_),
    .B1(_07449_),
    .B2(_06507_),
    .C1(_07451_),
    .C2(_07452_),
    .ZN(_07453_));
 MUX2_X1 _16712_ (.A(_07443_),
    .B(_07453_),
    .S(_06540_),
    .Z(_07454_));
 CLKBUF_X3 _16713_ (.A(_06572_),
    .Z(_07455_));
 MUX2_X1 _16714_ (.A(_07431_),
    .B(_07454_),
    .S(_07455_),
    .Z(_07456_));
 BUF_X4 _16715_ (.A(_06551_),
    .Z(_07457_));
 NAND2_X1 _16716_ (.A1(_07416_),
    .A2(_07457_),
    .ZN(_07458_));
 CLKBUF_X3 _16717_ (.A(_06524_),
    .Z(_07459_));
 BUF_X4 _16718_ (.A(_07459_),
    .Z(_07460_));
 MUX2_X1 _16719_ (.A(_07427_),
    .B(_07376_),
    .S(_06505_),
    .Z(_07461_));
 NOR2_X1 _16720_ (.A1(_07460_),
    .A2(_07461_),
    .ZN(_07462_));
 NAND2_X1 _16721_ (.A1(_14704_),
    .A2(_07379_),
    .ZN(_07463_));
 NAND2_X2 _16722_ (.A1(_06462_),
    .A2(_06505_),
    .ZN(_07464_));
 AND3_X1 _16723_ (.A1(_06525_),
    .A2(_07463_),
    .A3(_07464_),
    .ZN(_07465_));
 INV_X2 _16724_ (.A(_14694_),
    .ZN(_07466_));
 CLKBUF_X3 _16725_ (.A(_07378_),
    .Z(_07467_));
 NOR2_X1 _16726_ (.A1(_07466_),
    .A2(_07467_),
    .ZN(_07468_));
 OAI21_X1 _16727_ (.A(_07459_),
    .B1(_07412_),
    .B2(_07381_),
    .ZN(_07469_));
 OAI21_X1 _16728_ (.A(_07416_),
    .B1(_07468_),
    .B2(_07469_),
    .ZN(_07470_));
 BUF_X4 clone39 (.A(net600),
    .Z(net39));
 INV_X4 _16730_ (.A(_14701_),
    .ZN(_07472_));
 NAND2_X4 _16731_ (.A1(_06503_),
    .A2(_07410_),
    .ZN(_07473_));
 NOR2_X1 _16732_ (.A1(_07472_),
    .A2(_07473_),
    .ZN(_07474_));
 OAI33_X1 _16733_ (.A1(_07458_),
    .A2(_07462_),
    .A3(_07465_),
    .B1(_07470_),
    .B2(_07474_),
    .B3(_07457_),
    .ZN(_07475_));
 BUF_X8 _16734_ (.A(_06505_),
    .Z(_07476_));
 BUF_X4 _16735_ (.A(_07476_),
    .Z(_07477_));
 NOR3_X1 _16736_ (.A1(_14701_),
    .A2(_07389_),
    .A3(_07394_),
    .ZN(_07478_));
 AOI21_X2 _16737_ (.A(_14710_),
    .B1(_07384_),
    .B2(_07385_),
    .ZN(_07479_));
 OAI21_X1 _16738_ (.A(_07477_),
    .B1(_07478_),
    .B2(_07479_),
    .ZN(_07480_));
 AOI21_X1 _16739_ (.A(_07452_),
    .B1(_07419_),
    .B2(_07383_),
    .ZN(_07481_));
 AOI21_X1 _16740_ (.A(_07417_),
    .B1(_07480_),
    .B2(_07481_),
    .ZN(_07482_));
 BUF_X4 _16741_ (.A(_07410_),
    .Z(_07483_));
 BUF_X4 _16742_ (.A(_07483_),
    .Z(_07484_));
 INV_X2 _16743_ (.A(_14706_),
    .ZN(_07485_));
 AOI21_X1 _16744_ (.A(_07448_),
    .B1(_07484_),
    .B2(_07485_),
    .ZN(_07486_));
 BUF_X4 _16745_ (.A(_07378_),
    .Z(_07487_));
 CLKBUF_X3 _16746_ (.A(_07487_),
    .Z(_07488_));
 OAI221_X1 _16747_ (.A(_07452_),
    .B1(_07473_),
    .B2(net1238),
    .C1(_07486_),
    .C2(_07488_),
    .ZN(_07489_));
 AOI21_X1 _16748_ (.A(_07475_),
    .B1(_07482_),
    .B2(_07489_),
    .ZN(_07490_));
 CLKBUF_X3 _16749_ (.A(_07382_),
    .Z(_07491_));
 INV_X1 _16750_ (.A(_14710_),
    .ZN(_07492_));
 MUX2_X1 _16751_ (.A(_07492_),
    .B(net5),
    .S(_07378_),
    .Z(_07493_));
 NOR2_X1 _16752_ (.A1(_00385_),
    .A2(_07493_),
    .ZN(_07494_));
 INV_X1 _16753_ (.A(_07387_),
    .ZN(_07495_));
 NOR2_X1 _16754_ (.A1(_07495_),
    .A2(_06507_),
    .ZN(_07496_));
 CLKBUF_X3 _16755_ (.A(_07483_),
    .Z(_07497_));
 OAI21_X1 _16756_ (.A(_07497_),
    .B1(_07487_),
    .B2(_07377_),
    .ZN(_07498_));
 CLKBUF_X3 _16757_ (.A(_14696_),
    .Z(_07499_));
 CLKBUF_X3 _16758_ (.A(_07499_),
    .Z(_07500_));
 NOR2_X1 _16759_ (.A1(_07500_),
    .A2(_07487_),
    .ZN(_07501_));
 OAI22_X1 _16760_ (.A1(_07496_),
    .A2(_07498_),
    .B1(_07501_),
    .B2(_07469_),
    .ZN(_07502_));
 OAI221_X1 _16761_ (.A(_07491_),
    .B1(_07470_),
    .B2(_07494_),
    .C1(_07502_),
    .C2(_07417_),
    .ZN(_07503_));
 NOR2_X2 _16762_ (.A1(_06503_),
    .A2(_07410_),
    .ZN(_07504_));
 OAI22_X4 _16763_ (.A1(_06449_),
    .A2(net1054),
    .B1(_07388_),
    .B2(_07393_),
    .ZN(_07505_));
 NAND3_X2 _16764_ (.A1(_07387_),
    .A2(_06509_),
    .A3(_06521_),
    .ZN(_07506_));
 NAND2_X1 _16765_ (.A1(_07505_),
    .A2(_07506_),
    .ZN(_07507_));
 AOI221_X1 _16766_ (.A(_06538_),
    .B1(_07504_),
    .B2(_07472_),
    .C1(_07507_),
    .C2(_07467_),
    .ZN(_07508_));
 NAND3_X4 _16767_ (.A1(_07433_),
    .A2(_06509_),
    .A3(_06521_),
    .ZN(_07509_));
 AOI21_X1 _16768_ (.A(_07467_),
    .B1(_07505_),
    .B2(_07509_),
    .ZN(_07510_));
 OAI21_X1 _16769_ (.A(_07395_),
    .B1(_07497_),
    .B2(_07500_),
    .ZN(_07511_));
 AOI21_X1 _16770_ (.A(_07510_),
    .B1(_07511_),
    .B2(_07488_),
    .ZN(_07512_));
 AOI21_X1 _16771_ (.A(_07508_),
    .B1(_07512_),
    .B2(_06540_),
    .ZN(_07513_));
 OAI21_X1 _16772_ (.A(_07503_),
    .B1(_07513_),
    .B2(_07491_),
    .ZN(_07514_));
 MUX2_X1 _16773_ (.A(_07490_),
    .B(_07514_),
    .S(_07455_),
    .Z(_07515_));
 MUX2_X1 _16774_ (.A(_07456_),
    .B(_07515_),
    .S(_00388_),
    .Z(_00008_));
 INV_X2 _16775_ (.A(_06562_),
    .ZN(_07516_));
 NOR2_X1 _16776_ (.A1(_07516_),
    .A2(_00389_),
    .ZN(_07517_));
 CLKBUF_X3 _16777_ (.A(_07417_),
    .Z(_07518_));
 NAND3_X4 _16778_ (.A1(_14701_),
    .A2(_06509_),
    .A3(_06521_),
    .ZN(_07519_));
 NAND3_X1 _16779_ (.A1(_07412_),
    .A2(_07505_),
    .A3(_07519_),
    .ZN(_07520_));
 NAND2_X1 _16780_ (.A1(net14),
    .A2(_07460_),
    .ZN(_07521_));
 INV_X1 _16781_ (.A(_07383_),
    .ZN(_07522_));
 CLKBUF_X3 _16782_ (.A(_07497_),
    .Z(_07523_));
 NAND2_X1 _16783_ (.A1(_07522_),
    .A2(_07523_),
    .ZN(_07524_));
 NAND3_X1 _16784_ (.A1(_14712_),
    .A2(_07521_),
    .A3(_07524_),
    .ZN(_07525_));
 NAND4_X1 _16785_ (.A1(_07518_),
    .A2(_00387_),
    .A3(_07520_),
    .A4(_07525_),
    .ZN(_07526_));
 NOR3_X2 _16786_ (.A1(_06507_),
    .A2(_07402_),
    .A3(_07448_),
    .ZN(_07527_));
 AOI21_X1 _16787_ (.A(_07479_),
    .B1(_00385_),
    .B2(_07383_),
    .ZN(_07528_));
 AOI21_X1 _16788_ (.A(_07527_),
    .B1(_07528_),
    .B2(_14717_),
    .ZN(_07529_));
 NAND3_X2 _16789_ (.A1(_14694_),
    .A2(_07384_),
    .A3(_07385_),
    .ZN(_07530_));
 OAI21_X1 _16790_ (.A(_07530_),
    .B1(_07460_),
    .B2(_14710_),
    .ZN(_07531_));
 NAND3_X4 _16791_ (.A1(_07426_),
    .A2(_06509_),
    .A3(_06521_),
    .ZN(_07532_));
 OAI21_X1 _16792_ (.A(_07532_),
    .B1(_07460_),
    .B2(_07500_),
    .ZN(_07533_));
 BUF_X4 _16793_ (.A(_07477_),
    .Z(_07534_));
 MUX2_X1 _16794_ (.A(_07531_),
    .B(_07533_),
    .S(_07534_),
    .Z(_07535_));
 MUX2_X1 _16795_ (.A(_07529_),
    .B(_07535_),
    .S(_07491_),
    .Z(_07536_));
 OAI21_X1 _16796_ (.A(_07526_),
    .B1(_07536_),
    .B2(_07518_),
    .ZN(_07537_));
 CLKBUF_X3 _16797_ (.A(_07457_),
    .Z(_07538_));
 NOR2_X1 _16798_ (.A1(_06540_),
    .A2(_07538_),
    .ZN(_07539_));
 AOI21_X1 _16799_ (.A(_07466_),
    .B1(_07384_),
    .B2(_07385_),
    .ZN(_07540_));
 OAI21_X1 _16800_ (.A(_14717_),
    .B1(_07540_),
    .B2(_07448_),
    .ZN(_07541_));
 NAND3_X2 _16801_ (.A1(_14698_),
    .A2(_07487_),
    .A3(_07484_),
    .ZN(_07542_));
 AND3_X1 _16802_ (.A1(_07539_),
    .A2(_07541_),
    .A3(_07542_),
    .ZN(_07543_));
 OAI21_X1 _16803_ (.A(_07517_),
    .B1(_07537_),
    .B2(_07543_),
    .ZN(_07544_));
 NAND2_X2 _16804_ (.A1(_06538_),
    .A2(_06551_),
    .ZN(_07545_));
 AOI21_X1 _16805_ (.A(_07545_),
    .B1(_07405_),
    .B2(_07500_),
    .ZN(_07546_));
 MUX2_X1 _16806_ (.A(net32),
    .B(_14703_),
    .S(_00385_),
    .Z(_07547_));
 OAI21_X1 _16807_ (.A(_07546_),
    .B1(_07547_),
    .B2(_14712_),
    .ZN(_07548_));
 NOR2_X2 _16808_ (.A1(_07416_),
    .A2(_07457_),
    .ZN(_07549_));
 NOR2_X1 _16809_ (.A1(_14717_),
    .A2(_07402_),
    .ZN(_07550_));
 OAI21_X1 _16810_ (.A(_07550_),
    .B1(_07523_),
    .B2(net1238),
    .ZN(_07551_));
 OAI21_X2 _16811_ (.A(net955),
    .B1(_07389_),
    .B2(_07394_),
    .ZN(_07552_));
 NAND3_X1 _16812_ (.A1(_07444_),
    .A2(_07532_),
    .A3(_07552_),
    .ZN(_07553_));
 NAND3_X1 _16813_ (.A1(_07549_),
    .A2(_07551_),
    .A3(_07553_),
    .ZN(_07554_));
 NAND4_X1 _16814_ (.A1(_00388_),
    .A2(_00389_),
    .A3(_07548_),
    .A4(_07554_),
    .ZN(_07555_));
 NAND2_X4 _16815_ (.A1(_07378_),
    .A2(_07428_),
    .ZN(_07556_));
 AOI21_X1 _16816_ (.A(net1237),
    .B1(_07523_),
    .B2(net1238),
    .ZN(_07557_));
 OAI221_X1 _16817_ (.A(_00387_),
    .B1(_07556_),
    .B2(net32),
    .C1(_07557_),
    .C2(_14712_),
    .ZN(_07558_));
 XNOR2_X2 _16818_ (.A(_06505_),
    .B(_06524_),
    .ZN(_07559_));
 OAI22_X1 _16819_ (.A1(net1232),
    .A2(_07473_),
    .B1(_07559_),
    .B2(_14693_),
    .ZN(_07560_));
 NOR2_X1 _16820_ (.A1(net13),
    .A2(_07483_),
    .ZN(_07561_));
 AOI21_X1 _16821_ (.A(_07560_),
    .B1(_07561_),
    .B2(_14693_),
    .ZN(_07562_));
 OAI21_X1 _16822_ (.A(_07558_),
    .B1(_07562_),
    .B2(_00387_),
    .ZN(_07563_));
 AND2_X1 _16823_ (.A1(_07518_),
    .A2(_07563_),
    .ZN(_07564_));
 NAND2_X2 _16824_ (.A1(net1231),
    .A2(_07412_),
    .ZN(_07565_));
 NAND3_X1 _16825_ (.A1(_07523_),
    .A2(_07463_),
    .A3(_07565_),
    .ZN(_07566_));
 NOR3_X1 _16826_ (.A1(_14722_),
    .A2(_07497_),
    .A3(_07457_),
    .ZN(_07567_));
 NOR2_X1 _16827_ (.A1(_06540_),
    .A2(_07567_),
    .ZN(_07568_));
 NAND3_X1 _16828_ (.A1(_07412_),
    .A2(_07505_),
    .A3(_07530_),
    .ZN(_07569_));
 NAND3_X1 _16829_ (.A1(_07378_),
    .A2(_07506_),
    .A3(_07552_),
    .ZN(_07570_));
 AND2_X1 _16830_ (.A1(_07569_),
    .A2(_07570_),
    .ZN(_07571_));
 OAI21_X1 _16831_ (.A(_07520_),
    .B1(_07450_),
    .B2(_07444_),
    .ZN(_07572_));
 MUX2_X1 _16832_ (.A(_07571_),
    .B(_07572_),
    .S(_07382_),
    .Z(_07573_));
 AOI221_X2 _16833_ (.A(_06573_),
    .B1(_07566_),
    .B2(_07568_),
    .C1(_07573_),
    .C2(_00386_),
    .ZN(_07574_));
 NAND3_X1 _16834_ (.A1(_14693_),
    .A2(_14703_),
    .A3(_07497_),
    .ZN(_07575_));
 NOR3_X2 _16835_ (.A1(_07423_),
    .A2(_07389_),
    .A3(_07394_),
    .ZN(_07576_));
 AOI21_X1 _16836_ (.A(_07576_),
    .B1(_07497_),
    .B2(net13),
    .ZN(_07577_));
 OAI21_X1 _16837_ (.A(_07575_),
    .B1(_07577_),
    .B2(_07534_),
    .ZN(_07578_));
 OAI21_X2 _16838_ (.A(_07472_),
    .B1(_07389_),
    .B2(_07394_),
    .ZN(_07579_));
 AOI21_X2 _16839_ (.A(_06506_),
    .B1(_07509_),
    .B2(_07579_),
    .ZN(_07580_));
 AOI21_X1 _16840_ (.A(_07580_),
    .B1(_07511_),
    .B2(_07534_),
    .ZN(_07581_));
 MUX2_X1 _16841_ (.A(_07578_),
    .B(_07581_),
    .S(_07452_),
    .Z(_07582_));
 AND2_X1 _16842_ (.A1(_14713_),
    .A2(_06525_),
    .ZN(_07583_));
 MUX2_X1 _16843_ (.A(_07472_),
    .B(net13),
    .S(_07412_),
    .Z(_07584_));
 AOI21_X1 _16844_ (.A(_07583_),
    .B1(_07584_),
    .B2(_07484_),
    .ZN(_07585_));
 NAND3_X1 _16845_ (.A1(_06507_),
    .A2(_07509_),
    .A3(_07579_),
    .ZN(_07586_));
 NAND2_X1 _16846_ (.A1(_07403_),
    .A2(_07586_),
    .ZN(_07587_));
 MUX2_X1 _16847_ (.A(_07585_),
    .B(_07587_),
    .S(_06552_),
    .Z(_07588_));
 MUX2_X1 _16848_ (.A(_07582_),
    .B(_07588_),
    .S(_00386_),
    .Z(_07589_));
 AOI21_X2 _16849_ (.A(_07574_),
    .B1(_07589_),
    .B2(_00389_),
    .ZN(_07590_));
 OAI221_X2 _16850_ (.A(_07544_),
    .B1(_07555_),
    .B2(_07564_),
    .C1(_07590_),
    .C2(_00388_),
    .ZN(_00009_));
 NOR2_X2 _16851_ (.A1(_06540_),
    .A2(_07452_),
    .ZN(_07591_));
 NAND2_X4 _16852_ (.A1(_07509_),
    .A2(_07552_),
    .ZN(_07592_));
 OAI221_X1 _16853_ (.A(_07591_),
    .B1(_07592_),
    .B2(_14712_),
    .C1(_07556_),
    .C2(net1240),
    .ZN(_07593_));
 AND3_X1 _16854_ (.A1(_07516_),
    .A2(_00389_),
    .A3(_07593_),
    .ZN(_07594_));
 AOI22_X2 _16855_ (.A1(_14718_),
    .A2(_00385_),
    .B1(_07419_),
    .B2(_07423_),
    .ZN(_07595_));
 NAND2_X2 _16856_ (.A1(_07416_),
    .A2(_07382_),
    .ZN(_07596_));
 NAND2_X1 _16857_ (.A1(_14703_),
    .A2(_07444_),
    .ZN(_07597_));
 OAI21_X1 _16858_ (.A(_07597_),
    .B1(_07534_),
    .B2(_07423_),
    .ZN(_07598_));
 MUX2_X1 _16859_ (.A(_14715_),
    .B(_07598_),
    .S(_00385_),
    .Z(_07599_));
 NAND2_X2 _16860_ (.A1(_07476_),
    .A2(_06524_),
    .ZN(_07600_));
 NOR2_X1 _16861_ (.A1(_14698_),
    .A2(_07600_),
    .ZN(_07601_));
 AOI221_X1 _16862_ (.A(_07601_),
    .B1(_07419_),
    .B2(_14704_),
    .C1(net32),
    .C2(_07441_),
    .ZN(_07602_));
 MUX2_X1 _16863_ (.A(_07599_),
    .B(_07602_),
    .S(_00387_),
    .Z(_07603_));
 OAI221_X2 _16864_ (.A(_07594_),
    .B1(_07595_),
    .B2(_07596_),
    .C1(_07518_),
    .C2(_07603_),
    .ZN(_07604_));
 AOI21_X4 _16865_ (.A(_07433_),
    .B1(_07384_),
    .B2(_07385_),
    .ZN(_07605_));
 OAI21_X2 _16866_ (.A(_06506_),
    .B1(_07397_),
    .B2(_07605_),
    .ZN(_07606_));
 MUX2_X1 _16867_ (.A(_07492_),
    .B(net5),
    .S(_07483_),
    .Z(_07607_));
 OAI21_X1 _16868_ (.A(_07606_),
    .B1(_07607_),
    .B2(_14717_),
    .ZN(_07608_));
 NOR2_X1 _16869_ (.A1(_07491_),
    .A2(_07608_),
    .ZN(_07609_));
 AND3_X1 _16870_ (.A1(_07534_),
    .A2(_07579_),
    .A3(_07521_),
    .ZN(_07610_));
 OAI21_X1 _16871_ (.A(_07506_),
    .B1(_07460_),
    .B2(_07500_),
    .ZN(_07611_));
 NOR2_X1 _16872_ (.A1(_14717_),
    .A2(_07611_),
    .ZN(_07612_));
 NOR3_X1 _16873_ (.A1(_00387_),
    .A2(_07610_),
    .A3(_07612_),
    .ZN(_07613_));
 NOR3_X1 _16874_ (.A1(_07518_),
    .A2(_07609_),
    .A3(_07613_),
    .ZN(_07614_));
 AOI21_X1 _16875_ (.A(_14717_),
    .B1(_07395_),
    .B2(_07530_),
    .ZN(_07615_));
 NOR2_X1 _16876_ (.A1(_07500_),
    .A2(_07600_),
    .ZN(_07616_));
 MUX2_X1 _16877_ (.A(_14701_),
    .B(_07495_),
    .S(_07476_),
    .Z(_07617_));
 OAI21_X1 _16878_ (.A(_07416_),
    .B1(_07617_),
    .B2(_07484_),
    .ZN(_07618_));
 OAI33_X1 _16879_ (.A1(_07458_),
    .A2(_07615_),
    .A3(_07616_),
    .B1(_07618_),
    .B2(_07462_),
    .B3(_00387_),
    .ZN(_07619_));
 NOR2_X1 _16880_ (.A1(_07614_),
    .A2(_07619_),
    .ZN(_07620_));
 NAND2_X1 _16881_ (.A1(_07516_),
    .A2(_07455_),
    .ZN(_07621_));
 NOR2_X1 _16882_ (.A1(_07485_),
    .A2(_07459_),
    .ZN(_07622_));
 MUX2_X1 _16883_ (.A(net4),
    .B(net5),
    .S(_07415_),
    .Z(_07623_));
 AOI211_X2 _16884_ (.A(_07487_),
    .B(_07622_),
    .C1(_07623_),
    .C2(_07460_),
    .ZN(_07624_));
 AND3_X1 _16885_ (.A1(_07500_),
    .A2(_07497_),
    .A3(_06539_),
    .ZN(_07625_));
 AOI21_X1 _16886_ (.A(net1240),
    .B1(_07484_),
    .B2(_06539_),
    .ZN(_07626_));
 NOR3_X1 _16887_ (.A1(_14717_),
    .A2(_07625_),
    .A3(_07626_),
    .ZN(_07627_));
 OAI21_X1 _16888_ (.A(_07491_),
    .B1(_07624_),
    .B2(_07627_),
    .ZN(_07628_));
 AOI21_X1 _16889_ (.A(_07402_),
    .B1(_07459_),
    .B2(_07485_),
    .ZN(_07629_));
 AOI21_X4 _16890_ (.A(_07499_),
    .B1(_06509_),
    .B2(_06521_),
    .ZN(_07630_));
 AOI21_X1 _16891_ (.A(_07630_),
    .B1(_06525_),
    .B2(net13),
    .ZN(_07631_));
 MUX2_X1 _16892_ (.A(_07629_),
    .B(_07631_),
    .S(_07467_),
    .Z(_07632_));
 OAI21_X1 _16893_ (.A(_07532_),
    .B1(_07460_),
    .B2(_07407_),
    .ZN(_07633_));
 AOI21_X1 _16894_ (.A(_07510_),
    .B1(_07633_),
    .B2(_07380_),
    .ZN(_07634_));
 MUX2_X1 _16895_ (.A(_07632_),
    .B(_07634_),
    .S(_07417_),
    .Z(_07635_));
 OAI21_X1 _16896_ (.A(_07628_),
    .B1(_07635_),
    .B2(_07491_),
    .ZN(_07636_));
 MUX2_X1 _16897_ (.A(_06462_),
    .B(_06505_),
    .S(_07376_),
    .Z(_07637_));
 MUX2_X1 _16898_ (.A(_14722_),
    .B(_07637_),
    .S(_07459_),
    .Z(_07638_));
 NAND2_X1 _16899_ (.A1(_07433_),
    .A2(_07379_),
    .ZN(_07639_));
 AOI21_X1 _16900_ (.A(_07483_),
    .B1(_07412_),
    .B2(_07423_),
    .ZN(_07640_));
 AOI22_X1 _16901_ (.A1(_14720_),
    .A2(_07497_),
    .B1(_07639_),
    .B2(_07640_),
    .ZN(_07641_));
 MUX2_X1 _16902_ (.A(_07638_),
    .B(_07641_),
    .S(_07457_),
    .Z(_07642_));
 OAI21_X1 _16903_ (.A(_07432_),
    .B1(_07428_),
    .B2(_07376_),
    .ZN(_07643_));
 MUX2_X1 _16904_ (.A(_07643_),
    .B(_07592_),
    .S(_07379_),
    .Z(_07644_));
 AOI21_X2 _16905_ (.A(_14715_),
    .B1(_06461_),
    .B2(_07476_),
    .ZN(_07645_));
 MUX2_X1 _16906_ (.A(_07461_),
    .B(_07645_),
    .S(_07459_),
    .Z(_07646_));
 MUX2_X1 _16907_ (.A(_07644_),
    .B(_07646_),
    .S(_07457_),
    .Z(_07647_));
 MUX2_X1 _16908_ (.A(_07642_),
    .B(_07647_),
    .S(_00386_),
    .Z(_07648_));
 MUX2_X1 _16909_ (.A(_07636_),
    .B(_07648_),
    .S(_00389_),
    .Z(_07649_));
 OAI221_X2 _16910_ (.A(_07604_),
    .B1(_07620_),
    .B2(_07621_),
    .C1(_07649_),
    .C2(_07516_),
    .ZN(_00010_));
 MUX2_X1 _16911_ (.A(net5),
    .B(_07476_),
    .S(net4),
    .Z(_07650_));
 AOI221_X1 _16912_ (.A(_06551_),
    .B1(_07405_),
    .B2(_07423_),
    .C1(_07650_),
    .C2(_07447_),
    .ZN(_07651_));
 AOI21_X1 _16913_ (.A(_07467_),
    .B1(_07432_),
    .B2(_07437_),
    .ZN(_07652_));
 NOR3_X1 _16914_ (.A1(_07444_),
    .A2(_07576_),
    .A3(_07605_),
    .ZN(_07653_));
 NOR3_X2 _16915_ (.A1(_07452_),
    .A2(_07652_),
    .A3(_07653_),
    .ZN(_07654_));
 OAI21_X1 _16916_ (.A(_07417_),
    .B1(_07651_),
    .B2(_07654_),
    .ZN(_07655_));
 NAND3_X1 _16917_ (.A1(_07499_),
    .A2(_07384_),
    .A3(_07385_),
    .ZN(_07656_));
 OAI21_X1 _16918_ (.A(_07407_),
    .B1(_07389_),
    .B2(_07394_),
    .ZN(_07657_));
 AOI21_X1 _16919_ (.A(_06506_),
    .B1(_07656_),
    .B2(_07657_),
    .ZN(_07658_));
 OAI21_X2 _16920_ (.A(_07434_),
    .B1(_07410_),
    .B2(_06476_),
    .ZN(_07659_));
 AOI21_X1 _16921_ (.A(_07658_),
    .B1(_07659_),
    .B2(_06507_),
    .ZN(_07660_));
 NAND2_X1 _16922_ (.A1(_06477_),
    .A2(_07428_),
    .ZN(_07661_));
 OAI221_X1 _16923_ (.A(_07606_),
    .B1(_07661_),
    .B2(net3),
    .C1(_07421_),
    .C2(_07473_),
    .ZN(_07662_));
 MUX2_X1 _16924_ (.A(_07660_),
    .B(_07662_),
    .S(_06552_),
    .Z(_07663_));
 OAI21_X1 _16925_ (.A(_07655_),
    .B1(_07663_),
    .B2(_07518_),
    .ZN(_07664_));
 OAI21_X4 _16926_ (.A(net1051),
    .B1(_07410_),
    .B2(net1224),
    .ZN(_07665_));
 AOI221_X2 _16927_ (.A(_07379_),
    .B1(_07665_),
    .B2(_06551_),
    .C1(_07445_),
    .C2(_06463_),
    .ZN(_07666_));
 AOI21_X1 _16928_ (.A(_07630_),
    .B1(_07397_),
    .B2(_06551_),
    .ZN(_07667_));
 AND2_X1 _16929_ (.A1(_07380_),
    .A2(_07667_),
    .ZN(_07668_));
 NOR3_X2 _16930_ (.A1(_07417_),
    .A2(_07666_),
    .A3(_07668_),
    .ZN(_07669_));
 OAI21_X1 _16931_ (.A(_07477_),
    .B1(_07397_),
    .B2(_07540_),
    .ZN(_07670_));
 NAND3_X2 _16932_ (.A1(_07385_),
    .A2(_07384_),
    .A3(_14706_),
    .ZN(_07671_));
 OAI21_X1 _16933_ (.A(_07671_),
    .B1(_07459_),
    .B2(_14704_),
    .ZN(_07672_));
 OAI21_X1 _16934_ (.A(_07670_),
    .B1(_07672_),
    .B2(_06507_),
    .ZN(_07673_));
 OAI21_X1 _16935_ (.A(_07412_),
    .B1(_07428_),
    .B2(_07376_),
    .ZN(_07674_));
 AOI222_X2 _16936_ (.A1(_07522_),
    .A2(_07504_),
    .B1(_07674_),
    .B2(net3),
    .C1(_07377_),
    .C2(_07419_),
    .ZN(_07675_));
 MUX2_X1 _16937_ (.A(_07673_),
    .B(_07675_),
    .S(_06552_),
    .Z(_07676_));
 AOI21_X1 _16938_ (.A(_07669_),
    .B1(_07676_),
    .B2(_07518_),
    .ZN(_07677_));
 MUX2_X1 _16939_ (.A(_07664_),
    .B(_07677_),
    .S(_07455_),
    .Z(_07678_));
 AOI221_X1 _16940_ (.A(_06551_),
    .B1(_07405_),
    .B2(net1232),
    .C1(_07645_),
    .C2(_07447_),
    .ZN(_07679_));
 MUX2_X1 _16941_ (.A(_07421_),
    .B(_07522_),
    .S(_07428_),
    .Z(_07680_));
 OAI21_X1 _16942_ (.A(_07509_),
    .B1(_06525_),
    .B2(_06463_),
    .ZN(_07681_));
 MUX2_X1 _16943_ (.A(_07680_),
    .B(_07681_),
    .S(_07487_),
    .Z(_07682_));
 AOI21_X1 _16944_ (.A(_07679_),
    .B1(_07682_),
    .B2(_07538_),
    .ZN(_07683_));
 NOR3_X1 _16945_ (.A1(_06461_),
    .A2(net1226),
    .A3(_06524_),
    .ZN(_07684_));
 MUX2_X1 _16946_ (.A(_06461_),
    .B(net1225),
    .S(_06523_),
    .Z(_07685_));
 AOI221_X1 _16947_ (.A(_07684_),
    .B1(_07685_),
    .B2(_07378_),
    .C1(_07504_),
    .C2(net12),
    .ZN(_07686_));
 NAND3_X2 _16948_ (.A1(_07477_),
    .A2(net1053),
    .A3(_07656_),
    .ZN(_07687_));
 OAI21_X1 _16949_ (.A(_07519_),
    .B1(_06525_),
    .B2(_06477_),
    .ZN(_07688_));
 OAI21_X2 _16950_ (.A(_07687_),
    .B1(_07688_),
    .B2(_07444_),
    .ZN(_07689_));
 MUX2_X1 _16951_ (.A(_07686_),
    .B(_07689_),
    .S(_06552_),
    .Z(_07690_));
 MUX2_X1 _16952_ (.A(_07683_),
    .B(_07690_),
    .S(_07417_),
    .Z(_07691_));
 NOR2_X2 _16953_ (.A1(_06503_),
    .A2(_06523_),
    .ZN(_07692_));
 AOI22_X1 _16954_ (.A1(_07407_),
    .A2(_07559_),
    .B1(_07692_),
    .B2(_14693_),
    .ZN(_07693_));
 AOI21_X1 _16955_ (.A(_07402_),
    .B1(_06507_),
    .B2(_14693_),
    .ZN(_07694_));
 OAI221_X1 _16956_ (.A(_07542_),
    .B1(_07694_),
    .B2(net12),
    .C1(_14698_),
    .C2(_07600_),
    .ZN(_07695_));
 AOI21_X1 _16957_ (.A(_07397_),
    .B1(_07380_),
    .B2(_14698_),
    .ZN(_07696_));
 OAI21_X1 _16958_ (.A(_07452_),
    .B1(_07696_),
    .B2(_07500_),
    .ZN(_07697_));
 OAI22_X1 _16959_ (.A1(_07491_),
    .A2(_07693_),
    .B1(_07695_),
    .B2(_07697_),
    .ZN(_07698_));
 NOR2_X1 _16960_ (.A1(_00386_),
    .A2(_07698_),
    .ZN(_07699_));
 AOI21_X1 _16961_ (.A(_14704_),
    .B1(_07384_),
    .B2(_07385_),
    .ZN(_07700_));
 NOR3_X2 _16962_ (.A1(_07444_),
    .A2(_07448_),
    .A3(_07700_),
    .ZN(_07701_));
 AOI21_X1 _16963_ (.A(_07701_),
    .B1(_07607_),
    .B2(_07534_),
    .ZN(_07702_));
 AOI21_X1 _16964_ (.A(_07380_),
    .B1(_07422_),
    .B2(_07434_),
    .ZN(_07703_));
 MUX2_X1 _16965_ (.A(_07702_),
    .B(_07703_),
    .S(_06552_),
    .Z(_07704_));
 OAI21_X1 _16966_ (.A(_07455_),
    .B1(_07704_),
    .B2(_07518_),
    .ZN(_07705_));
 OAI22_X1 _16967_ (.A1(_07455_),
    .A2(_07691_),
    .B1(_07699_),
    .B2(_07705_),
    .ZN(_07706_));
 MUX2_X1 _16968_ (.A(_07678_),
    .B(_07706_),
    .S(_07516_),
    .Z(_00011_));
 AOI21_X1 _16969_ (.A(_07483_),
    .B1(_07379_),
    .B2(_06463_),
    .ZN(_07707_));
 AOI21_X2 _16970_ (.A(_06538_),
    .B1(_07565_),
    .B2(_07707_),
    .ZN(_07708_));
 NOR2_X1 _16971_ (.A1(net12),
    .A2(_07444_),
    .ZN(_07709_));
 NOR2_X1 _16972_ (.A1(net1240),
    .A2(_07487_),
    .ZN(_07710_));
 OAI21_X1 _16973_ (.A(_07523_),
    .B1(_07709_),
    .B2(_07710_),
    .ZN(_07711_));
 NOR2_X1 _16974_ (.A1(_07534_),
    .A2(_07416_),
    .ZN(_07712_));
 AOI221_X2 _16975_ (.A(_06573_),
    .B1(_07708_),
    .B2(_07711_),
    .C1(_07712_),
    .C2(_07531_),
    .ZN(_07713_));
 AOI221_X2 _16976_ (.A(_06539_),
    .B1(_07477_),
    .B2(net3),
    .C1(_14724_),
    .C2(_07460_),
    .ZN(_07714_));
 OAI21_X1 _16977_ (.A(_07714_),
    .B1(_07473_),
    .B2(_07383_),
    .ZN(_07715_));
 OAI221_X1 _16978_ (.A(_00386_),
    .B1(_07479_),
    .B2(_07488_),
    .C1(_07523_),
    .C2(_07485_),
    .ZN(_07716_));
 NAND3_X1 _16979_ (.A1(_06573_),
    .A2(_07715_),
    .A3(_07716_),
    .ZN(_07717_));
 NAND2_X1 _16980_ (.A1(_00387_),
    .A2(_07717_),
    .ZN(_07718_));
 AOI221_X1 _16981_ (.A(_07416_),
    .B1(_07405_),
    .B2(_07383_),
    .C1(_14703_),
    .C2(_06507_),
    .ZN(_07719_));
 NOR2_X1 _16982_ (.A1(_14693_),
    .A2(_07523_),
    .ZN(_07720_));
 NAND2_X1 _16983_ (.A1(net14),
    .A2(_07488_),
    .ZN(_07721_));
 AOI21_X1 _16984_ (.A(_00386_),
    .B1(_07720_),
    .B2(_07721_),
    .ZN(_07722_));
 NOR2_X1 _16985_ (.A1(_14698_),
    .A2(_07488_),
    .ZN(_07723_));
 OAI21_X1 _16986_ (.A(net14),
    .B1(_07419_),
    .B2(_07723_),
    .ZN(_07724_));
 AOI21_X1 _16987_ (.A(_07719_),
    .B1(_07722_),
    .B2(_07724_),
    .ZN(_07725_));
 AOI221_X2 _16988_ (.A(_14698_),
    .B1(_14703_),
    .B2(_07380_),
    .C1(_07384_),
    .C2(_07385_),
    .ZN(_07726_));
 NOR3_X1 _16989_ (.A1(_07455_),
    .A2(_07725_),
    .A3(_07726_),
    .ZN(_07727_));
 NAND2_X1 _16990_ (.A1(_07476_),
    .A2(_07410_),
    .ZN(_07728_));
 OAI221_X1 _16991_ (.A(_07417_),
    .B1(_07728_),
    .B2(_14693_),
    .C1(_07630_),
    .C2(_14717_),
    .ZN(_07729_));
 OAI21_X1 _16992_ (.A(_07519_),
    .B1(_00385_),
    .B2(_07383_),
    .ZN(_07730_));
 MUX2_X1 _16993_ (.A(_07450_),
    .B(_07730_),
    .S(_07534_),
    .Z(_07731_));
 OAI21_X1 _16994_ (.A(_07729_),
    .B1(_07731_),
    .B2(_07518_),
    .ZN(_07732_));
 OAI21_X1 _16995_ (.A(_07491_),
    .B1(_00389_),
    .B2(_07732_),
    .ZN(_07733_));
 OAI221_X1 _16996_ (.A(_00388_),
    .B1(_07713_),
    .B2(_07718_),
    .C1(_07727_),
    .C2(_07733_),
    .ZN(_07734_));
 AND3_X1 _16997_ (.A1(_07444_),
    .A2(_07506_),
    .A3(_07579_),
    .ZN(_07735_));
 AOI21_X2 _16998_ (.A(_07630_),
    .B1(_00385_),
    .B2(_14703_),
    .ZN(_07736_));
 AOI21_X1 _16999_ (.A(_07735_),
    .B1(_07736_),
    .B2(_07488_),
    .ZN(_07737_));
 OAI21_X1 _17000_ (.A(_07538_),
    .B1(_14712_),
    .B2(_07407_),
    .ZN(_07738_));
 OAI221_X1 _17001_ (.A(_00386_),
    .B1(_00387_),
    .B2(_07737_),
    .C1(_07738_),
    .C2(_07580_),
    .ZN(_07739_));
 MUX2_X1 _17002_ (.A(_07611_),
    .B(_07665_),
    .S(_07488_),
    .Z(_07740_));
 MUX2_X1 _17003_ (.A(net1238),
    .B(net14),
    .S(_07460_),
    .Z(_07741_));
 AOI21_X1 _17004_ (.A(_07596_),
    .B1(_07741_),
    .B2(_14712_),
    .ZN(_07742_));
 AOI22_X2 _17005_ (.A1(_07740_),
    .A2(_07591_),
    .B1(_07742_),
    .B2(_07396_),
    .ZN(_07743_));
 AND2_X4 _17006_ (.A1(_07739_),
    .A2(_07743_),
    .ZN(_07744_));
 NAND2_X1 _17007_ (.A1(_07407_),
    .A2(_07405_),
    .ZN(_07745_));
 NAND3_X1 _17008_ (.A1(_07534_),
    .A2(_07538_),
    .A3(_07395_),
    .ZN(_07746_));
 OAI21_X1 _17009_ (.A(_07746_),
    .B1(_07397_),
    .B2(_07538_),
    .ZN(_07747_));
 AOI21_X1 _17010_ (.A(_07488_),
    .B1(_00385_),
    .B2(_07538_),
    .ZN(_07748_));
 AOI21_X1 _17011_ (.A(_14712_),
    .B1(_07445_),
    .B2(net14),
    .ZN(_07749_));
 OAI221_X1 _17012_ (.A(_07747_),
    .B1(_07748_),
    .B2(net14),
    .C1(_07749_),
    .C2(_14693_),
    .ZN(_07750_));
 AOI21_X1 _17013_ (.A(_07518_),
    .B1(_07745_),
    .B2(_07750_),
    .ZN(_07751_));
 NAND2_X1 _17014_ (.A1(_07437_),
    .A2(_07591_),
    .ZN(_07752_));
 NOR2_X1 _17015_ (.A1(net1232),
    .A2(_07556_),
    .ZN(_07753_));
 NOR2_X1 _17016_ (.A1(_14710_),
    .A2(_07728_),
    .ZN(_07754_));
 AOI21_X1 _17017_ (.A(_07397_),
    .B1(_07523_),
    .B2(_07383_),
    .ZN(_07755_));
 OAI221_X1 _17018_ (.A(_07539_),
    .B1(_07755_),
    .B2(_14717_),
    .C1(_07521_),
    .C2(_14693_),
    .ZN(_07756_));
 OAI221_X1 _17019_ (.A(_07455_),
    .B1(_07752_),
    .B2(_07753_),
    .C1(_07754_),
    .C2(_07756_),
    .ZN(_07757_));
 OAI22_X4 _17020_ (.A1(_07455_),
    .A2(_07744_),
    .B1(_07751_),
    .B2(_07757_),
    .ZN(_07758_));
 OAI21_X4 _17021_ (.A(_07734_),
    .B1(_00388_),
    .B2(_07758_),
    .ZN(_00012_));
 NAND2_X1 _17022_ (.A1(_07409_),
    .A2(_07532_),
    .ZN(_07759_));
 AOI221_X1 _17023_ (.A(_07415_),
    .B1(_07692_),
    .B2(_06477_),
    .C1(_07759_),
    .C2(_07378_),
    .ZN(_07760_));
 MUX2_X1 _17024_ (.A(_07499_),
    .B(_07522_),
    .S(_07428_),
    .Z(_07761_));
 AOI21_X1 _17025_ (.A(_07440_),
    .B1(_07761_),
    .B2(_07380_),
    .ZN(_07762_));
 AOI21_X1 _17026_ (.A(_07760_),
    .B1(_07762_),
    .B2(_07417_),
    .ZN(_07763_));
 NOR2_X1 _17027_ (.A1(_07497_),
    .A2(_06539_),
    .ZN(_07764_));
 NOR3_X1 _17028_ (.A1(_06463_),
    .A2(_07459_),
    .A3(_07415_),
    .ZN(_07765_));
 OAI21_X1 _17029_ (.A(net15),
    .B1(_07764_),
    .B2(_07765_),
    .ZN(_07766_));
 NAND4_X1 _17030_ (.A1(_14703_),
    .A2(_07487_),
    .A3(_07497_),
    .A4(_07416_),
    .ZN(_07767_));
 NOR2_X1 _17031_ (.A1(_06477_),
    .A2(_06538_),
    .ZN(_07768_));
 OAI21_X1 _17032_ (.A(_14698_),
    .B1(_07419_),
    .B2(_07768_),
    .ZN(_07769_));
 NOR2_X1 _17033_ (.A1(_07483_),
    .A2(_07415_),
    .ZN(_07770_));
 NAND3_X1 _17034_ (.A1(_07463_),
    .A2(_07565_),
    .A3(_07770_),
    .ZN(_07771_));
 NAND4_X1 _17035_ (.A1(_07766_),
    .A2(_07767_),
    .A3(_07769_),
    .A4(_07771_),
    .ZN(_07772_));
 MUX2_X1 _17036_ (.A(_07763_),
    .B(_07772_),
    .S(_07538_),
    .Z(_07773_));
 NAND3_X1 _17037_ (.A1(_07423_),
    .A2(_07467_),
    .A3(_07447_),
    .ZN(_07774_));
 NAND3_X1 _17038_ (.A1(_07457_),
    .A2(_07774_),
    .A3(_07670_),
    .ZN(_07775_));
 OAI21_X1 _17039_ (.A(_07432_),
    .B1(_07565_),
    .B2(_07460_),
    .ZN(_07776_));
 OAI21_X1 _17040_ (.A(_07775_),
    .B1(_07776_),
    .B2(_06552_),
    .ZN(_07777_));
 NOR3_X1 _17041_ (.A1(_07421_),
    .A2(_07388_),
    .A3(_07393_),
    .ZN(_07778_));
 NOR3_X1 _17042_ (.A1(_07476_),
    .A2(_07778_),
    .A3(_07630_),
    .ZN(_07779_));
 AOI21_X1 _17043_ (.A(_07467_),
    .B1(net1052),
    .B2(_07532_),
    .ZN(_07780_));
 OAI21_X1 _17044_ (.A(_07382_),
    .B1(_07780_),
    .B2(_07779_),
    .ZN(_07781_));
 OAI21_X1 _17045_ (.A(_07447_),
    .B1(_07477_),
    .B2(_07472_),
    .ZN(_07782_));
 OAI21_X1 _17046_ (.A(_07782_),
    .B1(_07556_),
    .B2(_07500_),
    .ZN(_07783_));
 OAI21_X1 _17047_ (.A(_07781_),
    .B1(_07783_),
    .B2(_07452_),
    .ZN(_07784_));
 MUX2_X1 _17048_ (.A(_07777_),
    .B(_07784_),
    .S(_06540_),
    .Z(_07785_));
 MUX2_X1 _17049_ (.A(_07773_),
    .B(_07785_),
    .S(_07455_),
    .Z(_07786_));
 OAI221_X1 _17050_ (.A(_07464_),
    .B1(_07394_),
    .B2(_07389_),
    .C1(net1241),
    .C2(_07477_),
    .ZN(_07787_));
 NAND2_X1 _17051_ (.A1(_07708_),
    .A2(_07787_),
    .ZN(_07788_));
 AOI21_X1 _17052_ (.A(_07779_),
    .B1(_07692_),
    .B2(_07466_),
    .ZN(_07789_));
 AOI21_X1 _17053_ (.A(_07457_),
    .B1(_07789_),
    .B2(_06539_),
    .ZN(_07790_));
 NAND3_X1 _17054_ (.A1(_07381_),
    .A2(_07477_),
    .A3(_07447_),
    .ZN(_07791_));
 OAI21_X1 _17055_ (.A(_06463_),
    .B1(_06477_),
    .B2(_07459_),
    .ZN(_07792_));
 AOI21_X1 _17056_ (.A(_06539_),
    .B1(_07791_),
    .B2(_07792_),
    .ZN(_07793_));
 OAI21_X1 _17057_ (.A(_07509_),
    .B1(_07428_),
    .B2(net5),
    .ZN(_07794_));
 OAI21_X1 _17058_ (.A(_07506_),
    .B1(_07428_),
    .B2(_07407_),
    .ZN(_07795_));
 MUX2_X1 _17059_ (.A(_07794_),
    .B(_07795_),
    .S(_07379_),
    .Z(_07796_));
 AOI21_X1 _17060_ (.A(_07793_),
    .B1(_07796_),
    .B2(_06540_),
    .ZN(_07797_));
 AOI221_X1 _17061_ (.A(_06573_),
    .B1(_07788_),
    .B2(_07790_),
    .C1(_07797_),
    .C2(_07538_),
    .ZN(_07798_));
 MUX2_X1 _17062_ (.A(_07499_),
    .B(_06477_),
    .S(_07483_),
    .Z(_07799_));
 OAI21_X1 _17063_ (.A(_07480_),
    .B1(_07799_),
    .B2(_06507_),
    .ZN(_07800_));
 MUX2_X1 _17064_ (.A(_07397_),
    .B(_07665_),
    .S(_06506_),
    .Z(_07801_));
 MUX2_X1 _17065_ (.A(_07800_),
    .B(_07801_),
    .S(_07452_),
    .Z(_07802_));
 AOI22_X1 _17066_ (.A1(net1238),
    .A2(_07484_),
    .B1(_07506_),
    .B2(_07467_),
    .ZN(_07803_));
 NOR2_X1 _17067_ (.A1(_06552_),
    .A2(_07803_),
    .ZN(_07804_));
 AND3_X1 _17068_ (.A1(_07467_),
    .A2(_07519_),
    .A3(_07657_),
    .ZN(_07805_));
 MUX2_X1 _17069_ (.A(_07423_),
    .B(_07381_),
    .S(_06525_),
    .Z(_07806_));
 AOI21_X1 _17070_ (.A(_07805_),
    .B1(_07806_),
    .B2(_07534_),
    .ZN(_07807_));
 AOI21_X1 _17071_ (.A(_07804_),
    .B1(_07807_),
    .B2(_07538_),
    .ZN(_07808_));
 MUX2_X1 _17072_ (.A(_07802_),
    .B(_07808_),
    .S(_00386_),
    .Z(_07809_));
 AOI21_X2 _17073_ (.A(_07798_),
    .B1(_07809_),
    .B2(_00389_),
    .ZN(_07810_));
 MUX2_X1 _17074_ (.A(_07786_),
    .B(_07810_),
    .S(_00388_),
    .Z(_00013_));
 OAI221_X1 _17075_ (.A(_06539_),
    .B1(_07600_),
    .B2(_07377_),
    .C1(_07672_),
    .C2(_07444_),
    .ZN(_07811_));
 AND3_X1 _17076_ (.A1(_07452_),
    .A2(_07618_),
    .A3(_07811_),
    .ZN(_07812_));
 MUX2_X1 _17077_ (.A(_07485_),
    .B(_06477_),
    .S(_06505_),
    .Z(_07813_));
 MUX2_X1 _17078_ (.A(_14714_),
    .B(_07813_),
    .S(_07447_),
    .Z(_07814_));
 OAI21_X1 _17079_ (.A(_07656_),
    .B1(_06525_),
    .B2(_14698_),
    .ZN(_07815_));
 AOI21_X1 _17080_ (.A(_07440_),
    .B1(_07815_),
    .B2(_07380_),
    .ZN(_07816_));
 MUX2_X1 _17081_ (.A(_07814_),
    .B(_07816_),
    .S(_06539_),
    .Z(_07817_));
 AOI21_X1 _17082_ (.A(_07812_),
    .B1(_07817_),
    .B2(_00387_),
    .ZN(_07818_));
 NAND3_X1 _17083_ (.A1(_07495_),
    .A2(_07476_),
    .A3(_07428_),
    .ZN(_07819_));
 OAI221_X1 _17084_ (.A(_07819_),
    .B1(_07559_),
    .B2(_07381_),
    .C1(net12),
    .C2(_07473_),
    .ZN(_07820_));
 MUX2_X1 _17085_ (.A(_07411_),
    .B(_07659_),
    .S(_07476_),
    .Z(_07821_));
 MUX2_X1 _17086_ (.A(_07820_),
    .B(_07821_),
    .S(_07457_),
    .Z(_07822_));
 MUX2_X1 _17087_ (.A(_07433_),
    .B(_07387_),
    .S(_07378_),
    .Z(_07823_));
 MUX2_X1 _17088_ (.A(_14718_),
    .B(_07823_),
    .S(_07447_),
    .Z(_07824_));
 OAI21_X1 _17089_ (.A(_07487_),
    .B1(_07561_),
    .B2(_07700_),
    .ZN(_07825_));
 AND2_X1 _17090_ (.A1(_07382_),
    .A2(_07819_),
    .ZN(_07826_));
 AOI22_X1 _17091_ (.A1(_06552_),
    .A2(_07824_),
    .B1(_07825_),
    .B2(_07826_),
    .ZN(_07827_));
 MUX2_X1 _17092_ (.A(_07822_),
    .B(_07827_),
    .S(_06540_),
    .Z(_07828_));
 MUX2_X1 _17093_ (.A(_07818_),
    .B(_07828_),
    .S(_06573_),
    .Z(_07829_));
 AOI22_X1 _17094_ (.A1(net1232),
    .A2(_07419_),
    .B1(_07441_),
    .B2(_14698_),
    .ZN(_07830_));
 NAND2_X1 _17095_ (.A1(_07407_),
    .A2(_07504_),
    .ZN(_07831_));
 NAND3_X1 _17096_ (.A1(_07549_),
    .A2(_07830_),
    .A3(_07831_),
    .ZN(_07832_));
 OAI21_X1 _17097_ (.A(_07671_),
    .B1(_07459_),
    .B2(_07383_),
    .ZN(_07833_));
 AOI221_X2 _17098_ (.A(_07545_),
    .B1(_07833_),
    .B2(_07477_),
    .C1(_07405_),
    .C2(_14710_),
    .ZN(_07834_));
 OR2_X1 _17099_ (.A1(_14703_),
    .A2(_07397_),
    .ZN(_07835_));
 OAI21_X1 _17100_ (.A(_07835_),
    .B1(_07556_),
    .B2(net14),
    .ZN(_07836_));
 AOI21_X1 _17101_ (.A(_07834_),
    .B1(_07836_),
    .B2(_07591_),
    .ZN(_07837_));
 MUX2_X1 _17102_ (.A(_07499_),
    .B(_07407_),
    .S(_07378_),
    .Z(_07838_));
 AOI21_X2 _17103_ (.A(_07596_),
    .B1(_07838_),
    .B2(_07484_),
    .ZN(_07839_));
 AOI21_X1 _17104_ (.A(_07523_),
    .B1(_07488_),
    .B2(net32),
    .ZN(_07840_));
 OAI21_X1 _17105_ (.A(_07840_),
    .B1(_14712_),
    .B2(_14710_),
    .ZN(_07841_));
 AOI21_X1 _17106_ (.A(_06572_),
    .B1(_07839_),
    .B2(_07841_),
    .ZN(_07842_));
 NAND3_X1 _17107_ (.A1(_07832_),
    .A2(_07837_),
    .A3(_07842_),
    .ZN(_07843_));
 AOI21_X1 _17108_ (.A(_06506_),
    .B1(_06525_),
    .B2(_06463_),
    .ZN(_07844_));
 AND2_X1 _17109_ (.A1(_06506_),
    .A2(_07665_),
    .ZN(_07845_));
 OAI22_X1 _17110_ (.A1(net3),
    .A2(_07661_),
    .B1(_07728_),
    .B2(_07499_),
    .ZN(_07846_));
 NOR2_X1 _17111_ (.A1(_06463_),
    .A2(_06506_),
    .ZN(_07847_));
 OAI33_X1 _17112_ (.A1(_07596_),
    .A2(_07844_),
    .A3(_07845_),
    .B1(_07846_),
    .B2(_07847_),
    .B3(_07545_),
    .ZN(_07848_));
 OAI221_X1 _17113_ (.A(_07464_),
    .B1(_07394_),
    .B2(_07389_),
    .C1(_07495_),
    .C2(_07477_),
    .ZN(_07849_));
 OAI21_X1 _17114_ (.A(_07849_),
    .B1(_07484_),
    .B2(_14713_),
    .ZN(_07850_));
 NOR2_X1 _17115_ (.A1(_14703_),
    .A2(_07844_),
    .ZN(_07851_));
 NOR2_X1 _17116_ (.A1(_07458_),
    .A2(_07851_),
    .ZN(_07852_));
 AOI21_X1 _17117_ (.A(_07601_),
    .B1(_07419_),
    .B2(_07423_),
    .ZN(_07853_));
 AOI221_X2 _17118_ (.A(_07848_),
    .B1(_07850_),
    .B2(_07549_),
    .C1(_07852_),
    .C2(_07853_),
    .ZN(_07854_));
 OAI21_X1 _17119_ (.A(_07843_),
    .B1(_07854_),
    .B2(_00389_),
    .ZN(_07855_));
 MUX2_X1 _17120_ (.A(_07829_),
    .B(_07855_),
    .S(_00388_),
    .Z(_00014_));
 OAI221_X1 _17121_ (.A(_07415_),
    .B1(_07473_),
    .B2(_07492_),
    .C1(net32),
    .C2(_07410_),
    .ZN(_07856_));
 OAI21_X1 _17122_ (.A(_07519_),
    .B1(_06524_),
    .B2(_07387_),
    .ZN(_07857_));
 MUX2_X1 _17123_ (.A(_07450_),
    .B(_07857_),
    .S(_06505_),
    .Z(_07858_));
 OAI21_X1 _17124_ (.A(_07856_),
    .B1(_07858_),
    .B2(_07415_),
    .ZN(_07859_));
 NAND2_X1 _17125_ (.A1(_06522_),
    .A2(_06538_),
    .ZN(_07860_));
 NAND2_X1 _17126_ (.A1(_06523_),
    .A2(_07415_),
    .ZN(_07861_));
 OAI21_X1 _17127_ (.A(_07860_),
    .B1(_07861_),
    .B2(net1226),
    .ZN(_07862_));
 NOR3_X1 _17128_ (.A1(_06505_),
    .A2(_06524_),
    .A3(_06538_),
    .ZN(_07863_));
 AOI221_X2 _17129_ (.A(_06573_),
    .B1(_07862_),
    .B2(net4),
    .C1(_07863_),
    .C2(_07466_),
    .ZN(_07864_));
 NAND3_X1 _17130_ (.A1(_07476_),
    .A2(_07483_),
    .A3(_07415_),
    .ZN(_07865_));
 AOI21_X1 _17131_ (.A(_06477_),
    .B1(_07556_),
    .B2(_07865_),
    .ZN(_07866_));
 NOR3_X1 _17132_ (.A1(_07447_),
    .A2(_07415_),
    .A3(_07464_),
    .ZN(_07867_));
 NOR2_X1 _17133_ (.A1(_07866_),
    .A2(_07867_),
    .ZN(_07868_));
 AOI221_X2 _17134_ (.A(_07382_),
    .B1(_06573_),
    .B2(_07859_),
    .C1(_07864_),
    .C2(_07868_),
    .ZN(_07869_));
 INV_X1 _17135_ (.A(_14720_),
    .ZN(_07870_));
 OAI21_X1 _17136_ (.A(_06539_),
    .B1(_00385_),
    .B2(_07870_),
    .ZN(_07871_));
 NOR3_X1 _17137_ (.A1(_07440_),
    .A2(_07527_),
    .A3(_07871_),
    .ZN(_07872_));
 OAI221_X1 _17138_ (.A(_07416_),
    .B1(_07394_),
    .B2(_07389_),
    .C1(_07485_),
    .C2(_07487_),
    .ZN(_07873_));
 OAI221_X1 _17139_ (.A(_06573_),
    .B1(_07709_),
    .B2(_07873_),
    .C1(_07861_),
    .C2(_14724_),
    .ZN(_07874_));
 AOI21_X1 _17140_ (.A(_07466_),
    .B1(_07473_),
    .B2(_07861_),
    .ZN(_07875_));
 AOI221_X2 _17141_ (.A(_07379_),
    .B1(_07483_),
    .B2(_07427_),
    .C1(_07770_),
    .C2(_07423_),
    .ZN(_07876_));
 OAI21_X1 _17142_ (.A(_06572_),
    .B1(_07712_),
    .B2(_07876_),
    .ZN(_07877_));
 OAI22_X1 _17143_ (.A1(_07872_),
    .A2(_07874_),
    .B1(_07875_),
    .B2(_07877_),
    .ZN(_07878_));
 AOI211_X2 _17144_ (.A(_07869_),
    .B(_00388_),
    .C1(_07878_),
    .C2(_07491_),
    .ZN(_07879_));
 NAND3_X1 _17145_ (.A1(_07380_),
    .A2(_07432_),
    .A3(_07437_),
    .ZN(_07880_));
 AND3_X1 _17146_ (.A1(_06552_),
    .A2(_07553_),
    .A3(_07880_),
    .ZN(_07881_));
 NOR2_X1 _17147_ (.A1(_07383_),
    .A2(_07380_),
    .ZN(_07882_));
 OAI21_X1 _17148_ (.A(_07409_),
    .B1(_07523_),
    .B2(net14),
    .ZN(_07883_));
 AOI21_X1 _17149_ (.A(_07882_),
    .B1(_07883_),
    .B2(_07488_),
    .ZN(_07884_));
 AOI21_X1 _17150_ (.A(_07881_),
    .B1(_07884_),
    .B2(_07491_),
    .ZN(_07885_));
 AOI21_X1 _17151_ (.A(_07447_),
    .B1(net13),
    .B2(net3),
    .ZN(_07886_));
 AOI22_X1 _17152_ (.A1(net1240),
    .A2(_07484_),
    .B1(_07597_),
    .B2(_07886_),
    .ZN(_07887_));
 MUX2_X1 _17153_ (.A(_06463_),
    .B(_06477_),
    .S(_07410_),
    .Z(_07888_));
 OAI21_X1 _17154_ (.A(_07671_),
    .B1(_06525_),
    .B2(_14694_),
    .ZN(_07889_));
 MUX2_X1 _17155_ (.A(_07888_),
    .B(_07889_),
    .S(_07467_),
    .Z(_07890_));
 MUX2_X1 _17156_ (.A(_07887_),
    .B(_07890_),
    .S(_07538_),
    .Z(_07891_));
 MUX2_X1 _17157_ (.A(_07885_),
    .B(_07891_),
    .S(_00386_),
    .Z(_07892_));
 OAI22_X2 _17158_ (.A1(_07407_),
    .A2(_07556_),
    .B1(_07736_),
    .B2(_14712_),
    .ZN(_07893_));
 AOI21_X1 _17159_ (.A(_07545_),
    .B1(_07550_),
    .B2(_07530_),
    .ZN(_07894_));
 AOI22_X2 _17160_ (.A1(_07591_),
    .A2(_07893_),
    .B1(_07894_),
    .B2(_07396_),
    .ZN(_07895_));
 OR2_X1 _17161_ (.A1(_07484_),
    .A2(_07645_),
    .ZN(_07896_));
 OAI221_X2 _17162_ (.A(_07542_),
    .B1(_07600_),
    .B2(_07500_),
    .C1(net12),
    .C2(_07559_),
    .ZN(_07897_));
 AOI221_X2 _17163_ (.A(_06573_),
    .B1(_07896_),
    .B2(_07839_),
    .C1(_07897_),
    .C2(_07549_),
    .ZN(_07898_));
 AOI22_X2 _17164_ (.A1(_00389_),
    .A2(_07892_),
    .B1(_07895_),
    .B2(_07898_),
    .ZN(_07899_));
 AOI21_X4 _17165_ (.A(_07879_),
    .B1(_07899_),
    .B2(_00388_),
    .ZN(_00015_));
 BUF_X8 _17166_ (.A(_06351_),
    .Z(_14726_));
 BUF_X16 _17167_ (.A(_06379_),
    .Z(_07900_));
 BUF_X16 _17168_ (.A(_07900_),
    .Z(_07901_));
 BUF_X16 _17169_ (.A(_07901_),
    .Z(_14746_));
 BUF_X8 _17170_ (.A(_06335_),
    .Z(_07902_));
 BUF_X4 rebuffer569 (.A(_15057_),
    .Z(net1032));
 BUF_X4 _17172_ (.A(_06411_),
    .Z(_07903_));
 BUF_X4 _17173_ (.A(_07903_),
    .Z(_07904_));
 BUF_X4 _17174_ (.A(_14729_),
    .Z(_07905_));
 INV_X8 _17175_ (.A(_07905_),
    .ZN(_07906_));
 BUF_X4 _17176_ (.A(_06398_),
    .Z(_07907_));
 NAND2_X2 _17177_ (.A1(_06381_),
    .A2(_07907_),
    .ZN(_07908_));
 NOR3_X1 _17178_ (.A1(_07906_),
    .A2(_06447_),
    .A3(_07908_),
    .ZN(_07909_));
 BUF_X4 _17179_ (.A(_06399_),
    .Z(_07910_));
 CLKBUF_X3 _17180_ (.A(_07910_),
    .Z(_07911_));
 AND3_X1 _17181_ (.A1(_14754_),
    .A2(_07911_),
    .A3(_06447_),
    .ZN(_07912_));
 BUF_X8 _17182_ (.A(_07905_),
    .Z(_07913_));
 NOR2_X4 _17183_ (.A1(_06218_),
    .A2(net116),
    .ZN(_07914_));
 BUF_X8 _17184_ (.A(_07914_),
    .Z(_07915_));
 BUF_X4 _17185_ (.A(_07915_),
    .Z(_07916_));
 NOR2_X1 _17186_ (.A1(net16),
    .A2(_06390_),
    .ZN(_07917_));
 NOR2_X1 _17187_ (.A1(_06245_),
    .A2(_06388_),
    .ZN(_07918_));
 MUX2_X2 _17188_ (.A(_07917_),
    .B(_07918_),
    .S(_06395_),
    .Z(_07919_));
 BUF_X8 _17189_ (.A(_07919_),
    .Z(_07920_));
 BUF_X4 _17190_ (.A(_07920_),
    .Z(_07921_));
 OAI221_X1 _17191_ (.A(_07913_),
    .B1(_07916_),
    .B2(_07921_),
    .C1(_06447_),
    .C2(_06351_),
    .ZN(_07922_));
 INV_X1 _17192_ (.A(net73),
    .ZN(_07923_));
 NAND2_X1 _17193_ (.A1(_06401_),
    .A2(_07923_),
    .ZN(_07924_));
 NAND2_X1 _17194_ (.A1(_06266_),
    .A2(_06344_),
    .ZN(_07925_));
 NAND2_X1 _17195_ (.A1(_06266_),
    .A2(_06342_),
    .ZN(_07926_));
 MUX2_X1 _17196_ (.A(_07925_),
    .B(_07926_),
    .S(_06349_),
    .Z(_07927_));
 AOI22_X4 _17197_ (.A1(_07924_),
    .A2(_07927_),
    .B1(_06385_),
    .B2(_06397_),
    .ZN(_07928_));
 OR3_X1 _17198_ (.A1(_07913_),
    .A2(_06446_),
    .A3(_07928_),
    .ZN(_07929_));
 AOI21_X1 _17199_ (.A(_06383_),
    .B1(_07922_),
    .B2(_07929_),
    .ZN(_07930_));
 NOR4_X2 _17200_ (.A1(_07904_),
    .A2(_07909_),
    .A3(_07912_),
    .A4(_07930_),
    .ZN(_07931_));
 BUF_X2 split101 (.A(_15306_),
    .Z(net101));
 OAI21_X2 _17202_ (.A(net1122),
    .B1(_07915_),
    .B2(_07920_),
    .ZN(_07933_));
 BUF_X4 _17203_ (.A(_06385_),
    .Z(_07934_));
 BUF_X4 _17204_ (.A(_06397_),
    .Z(_07935_));
 NAND3_X2 _17205_ (.A1(_14742_),
    .A2(_07934_),
    .A3(_07935_),
    .ZN(_07936_));
 NAND3_X2 _17206_ (.A1(_06381_),
    .A2(_07933_),
    .A3(_07936_),
    .ZN(_07937_));
 XNOR2_X1 _17207_ (.A(_14732_),
    .B(_00400_),
    .ZN(_07938_));
 OAI211_X2 _17208_ (.A(_06447_),
    .B(_07937_),
    .C1(_07938_),
    .C2(_14751_),
    .ZN(_07939_));
 BUF_X4 _17209_ (.A(_07913_),
    .Z(_07940_));
 NAND3_X1 _17210_ (.A1(_07940_),
    .A2(_06383_),
    .A3(_00400_),
    .ZN(_07941_));
 XNOR2_X2 _17211_ (.A(_06381_),
    .B(_06399_),
    .ZN(_07942_));
 CLKBUF_X3 _17212_ (.A(_14742_),
    .Z(_07943_));
 NAND2_X4 _17213_ (.A1(_07900_),
    .A2(_07907_),
    .ZN(_07944_));
 BUF_X4 clone27 (.A(net28),
    .Z(net27));
 OAI221_X1 _17215_ (.A(_07941_),
    .B1(_07942_),
    .B2(_07943_),
    .C1(_07944_),
    .C2(net99),
    .ZN(_07946_));
 OAI21_X1 _17216_ (.A(_07939_),
    .B1(_07946_),
    .B2(_06448_),
    .ZN(_07947_));
 CLKBUF_X3 _17217_ (.A(_07904_),
    .Z(_07948_));
 AOI21_X1 _17218_ (.A(_07931_),
    .B1(_07947_),
    .B2(_07948_),
    .ZN(_07949_));
 BUF_X4 _17219_ (.A(_07900_),
    .Z(_07950_));
 BUF_X2 split99 (.A(_14738_),
    .Z(net99));
 NOR3_X1 _17221_ (.A1(net1117),
    .A2(_07916_),
    .A3(_07921_),
    .ZN(_07952_));
 NOR3_X1 _17222_ (.A1(_07950_),
    .A2(_07928_),
    .A3(_07952_),
    .ZN(_07953_));
 OAI221_X1 _17223_ (.A(_06397_),
    .B1(_06334_),
    .B2(_06324_),
    .C1(_06267_),
    .C2(net116),
    .ZN(_07954_));
 CLKBUF_X3 _17224_ (.A(_07954_),
    .Z(_07955_));
 AND2_X1 _17225_ (.A1(_07933_),
    .A2(_07955_),
    .ZN(_07956_));
 CLKBUF_X3 _17226_ (.A(_06379_),
    .Z(_07957_));
 BUF_X4 _17227_ (.A(_07957_),
    .Z(_07958_));
 AOI21_X1 _17228_ (.A(_07953_),
    .B1(_07956_),
    .B2(_07958_),
    .ZN(_07959_));
 CLKBUF_X2 _17229_ (.A(_14728_),
    .Z(_07960_));
 CLKBUF_X3 _17230_ (.A(_07960_),
    .Z(_07961_));
 NAND2_X1 _17231_ (.A1(_07961_),
    .A2(_06382_),
    .ZN(_07962_));
 CLKBUF_X3 _17232_ (.A(_06379_),
    .Z(_07963_));
 AOI21_X1 _17233_ (.A(_07907_),
    .B1(_07963_),
    .B2(_06336_),
    .ZN(_07964_));
 AOI21_X2 _17234_ (.A(_06412_),
    .B1(_07962_),
    .B2(_07964_),
    .ZN(_07965_));
 BUF_X4 _17235_ (.A(_07907_),
    .Z(_07966_));
 BUF_X4 _17236_ (.A(_07966_),
    .Z(_07967_));
 CLKBUF_X3 _17237_ (.A(_14744_),
    .Z(_07968_));
 MUX2_X1 _17238_ (.A(_07968_),
    .B(_06352_),
    .S(_07900_),
    .Z(_07969_));
 NAND2_X1 _17239_ (.A1(_07967_),
    .A2(_07969_),
    .ZN(_07970_));
 AOI22_X1 _17240_ (.A1(_06414_),
    .A2(_07959_),
    .B1(_07965_),
    .B2(_07970_),
    .ZN(_07971_));
 INV_X1 _17241_ (.A(_07960_),
    .ZN(_07972_));
 BUF_X4 _17242_ (.A(_06381_),
    .Z(_07973_));
 BUF_X4 _17243_ (.A(_07973_),
    .Z(_07974_));
 BUF_X4 _17244_ (.A(_07907_),
    .Z(_07975_));
 NOR2_X1 _17245_ (.A1(_07975_),
    .A2(_06412_),
    .ZN(_07976_));
 NAND3_X1 _17246_ (.A1(_07972_),
    .A2(_07974_),
    .A3(_07976_),
    .ZN(_07977_));
 NOR3_X4 _17247_ (.A1(_07906_),
    .A2(_07915_),
    .A3(_07920_),
    .ZN(_07978_));
 NOR2_X1 _17248_ (.A1(_07957_),
    .A2(_06400_),
    .ZN(_07979_));
 BUF_X4 rebuffer748 (.A(_15131_),
    .Z(net1211));
 BUF_X4 _17250_ (.A(_14740_),
    .Z(_07981_));
 AOI21_X1 _17251_ (.A(_07978_),
    .B1(_07979_),
    .B2(_07981_),
    .ZN(_07982_));
 BUF_X8 _17252_ (.A(_14735_),
    .Z(_07983_));
 OAI21_X2 _17253_ (.A(net1163),
    .B1(_07916_),
    .B2(_07921_),
    .ZN(_07984_));
 OAI21_X1 _17254_ (.A(_07911_),
    .B1(_06412_),
    .B2(net39),
    .ZN(_07985_));
 AND2_X1 _17255_ (.A1(_07984_),
    .A2(_07985_),
    .ZN(_07986_));
 OAI221_X1 _17256_ (.A(_07977_),
    .B1(_07982_),
    .B2(_07904_),
    .C1(_14751_),
    .C2(_07986_),
    .ZN(_07987_));
 MUX2_X1 _17257_ (.A(_07971_),
    .B(_07987_),
    .S(_06447_),
    .Z(_07988_));
 MUX2_X1 _17258_ (.A(_07949_),
    .B(_07988_),
    .S(_00403_),
    .Z(_07989_));
 MUX2_X1 _17259_ (.A(_06351_),
    .B(_06379_),
    .S(net600),
    .Z(_07990_));
 XNOR2_X1 _17260_ (.A(_07975_),
    .B(_07990_),
    .ZN(_07991_));
 INV_X1 _17261_ (.A(net19),
    .ZN(_07992_));
 AOI221_X1 _17262_ (.A(_06334_),
    .B1(_06385_),
    .B2(_06397_),
    .C1(_07992_),
    .C2(_06401_),
    .ZN(_07993_));
 CLKBUF_X3 _17263_ (.A(_07993_),
    .Z(_07994_));
 OR2_X2 _17264_ (.A1(_07978_),
    .A2(_07994_),
    .ZN(_07995_));
 AOI21_X4 _17265_ (.A(_14733_),
    .B1(_06385_),
    .B2(_06397_),
    .ZN(_07996_));
 INV_X4 _17266_ (.A(net1169),
    .ZN(_07997_));
 NOR3_X4 _17267_ (.A1(_07997_),
    .A2(_07915_),
    .A3(_07920_),
    .ZN(_07998_));
 OR2_X2 _17268_ (.A1(_07996_),
    .A2(_07998_),
    .ZN(_07999_));
 MUX2_X1 _17269_ (.A(_07995_),
    .B(_07999_),
    .S(_07963_),
    .Z(_08000_));
 MUX2_X1 _17270_ (.A(_07991_),
    .B(_08000_),
    .S(_06438_),
    .Z(_08001_));
 NAND2_X4 _17271_ (.A1(_06381_),
    .A2(_06399_),
    .ZN(_08002_));
 INV_X2 _17272_ (.A(_14733_),
    .ZN(_08003_));
 NOR3_X4 _17273_ (.A1(_07914_),
    .A2(_08003_),
    .A3(_07919_),
    .ZN(_08004_));
 AOI21_X1 _17274_ (.A(_08004_),
    .B1(_07967_),
    .B2(_06336_),
    .ZN(_08005_));
 OAI221_X1 _17275_ (.A(_06438_),
    .B1(_08002_),
    .B2(net1163),
    .C1(_08005_),
    .C2(_06383_),
    .ZN(_08006_));
 BUF_X4 _17276_ (.A(_06380_),
    .Z(_08007_));
 BUF_X4 _17277_ (.A(_08007_),
    .Z(_08008_));
 NAND3_X4 _17278_ (.A1(_14738_),
    .A2(_07934_),
    .A3(_07935_),
    .ZN(_08009_));
 OAI21_X4 _17279_ (.A(_07906_),
    .B1(_07916_),
    .B2(_07921_),
    .ZN(_08010_));
 NAND3_X1 _17280_ (.A1(_08008_),
    .A2(_08009_),
    .A3(_08010_),
    .ZN(_08011_));
 OAI21_X2 _17281_ (.A(_07960_),
    .B1(_07915_),
    .B2(_07920_),
    .ZN(_08012_));
 NAND3_X1 _17282_ (.A1(_07950_),
    .A2(_07936_),
    .A3(_08012_),
    .ZN(_08013_));
 AND2_X1 _17283_ (.A1(_08011_),
    .A2(_08013_),
    .ZN(_08014_));
 OAI21_X1 _17284_ (.A(_08006_),
    .B1(_08014_),
    .B2(_06438_),
    .ZN(_08015_));
 MUX2_X1 _17285_ (.A(_08001_),
    .B(_08015_),
    .S(_07904_),
    .Z(_08016_));
 NAND3_X1 _17286_ (.A1(_07981_),
    .A2(_07963_),
    .A3(_06400_),
    .ZN(_08017_));
 AOI21_X2 _17287_ (.A(_14744_),
    .B1(_07934_),
    .B2(_07935_),
    .ZN(_08018_));
 OR2_X1 _17288_ (.A1(_08004_),
    .A2(_08018_),
    .ZN(_08019_));
 OAI21_X1 _17289_ (.A(_08017_),
    .B1(_08019_),
    .B2(_07950_),
    .ZN(_08020_));
 NOR4_X4 _17290_ (.A1(_06324_),
    .A2(net1016),
    .A3(_07914_),
    .A4(_07919_),
    .ZN(_08021_));
 OAI21_X1 _17291_ (.A(_08007_),
    .B1(_07928_),
    .B2(_08021_),
    .ZN(_08022_));
 OAI21_X2 _17292_ (.A(_07905_),
    .B1(_07915_),
    .B2(_07920_),
    .ZN(_08023_));
 NAND3_X1 _17293_ (.A1(_07957_),
    .A2(_08009_),
    .A3(_08023_),
    .ZN(_08024_));
 NAND2_X1 _17294_ (.A1(_08022_),
    .A2(_08024_),
    .ZN(_08025_));
 MUX2_X1 _17295_ (.A(_08020_),
    .B(_08025_),
    .S(_06438_),
    .Z(_08026_));
 AOI21_X1 _17296_ (.A(_07996_),
    .B1(_07910_),
    .B2(_07968_),
    .ZN(_08027_));
 OAI22_X1 _17297_ (.A1(_14738_),
    .A2(_07944_),
    .B1(_08027_),
    .B2(_07957_),
    .ZN(_08028_));
 NOR3_X4 _17298_ (.A1(_07983_),
    .A2(_07915_),
    .A3(_07920_),
    .ZN(_08029_));
 OAI21_X2 _17299_ (.A(_06382_),
    .B1(_08018_),
    .B2(_08029_),
    .ZN(_08030_));
 NAND3_X1 _17300_ (.A1(_07943_),
    .A2(_07963_),
    .A3(_07966_),
    .ZN(_08031_));
 AND2_X2 _17301_ (.A1(_08030_),
    .A2(_08031_),
    .ZN(_08032_));
 MUX2_X1 _17302_ (.A(_08028_),
    .B(_08032_),
    .S(_06438_),
    .Z(_08033_));
 BUF_X4 _17303_ (.A(_06413_),
    .Z(_08034_));
 MUX2_X1 _17304_ (.A(_08026_),
    .B(_08033_),
    .S(_08034_),
    .Z(_08035_));
 MUX2_X1 _17305_ (.A(_08016_),
    .B(_08035_),
    .S(_00404_),
    .Z(_08036_));
 MUX2_X1 _17306_ (.A(_07989_),
    .B(_08036_),
    .S(_00402_),
    .Z(_00016_));
 OR3_X1 _17307_ (.A1(_14756_),
    .A2(_07975_),
    .A3(_06426_),
    .ZN(_08037_));
 NAND2_X1 _17308_ (.A1(net99),
    .A2(_07950_),
    .ZN(_08038_));
 NAND3_X1 _17309_ (.A1(_07967_),
    .A2(_07962_),
    .A3(_08038_),
    .ZN(_08039_));
 AOI21_X1 _17310_ (.A(_06413_),
    .B1(_08037_),
    .B2(_08039_),
    .ZN(_08040_));
 NAND3_X1 _17311_ (.A1(net1122),
    .A2(_07934_),
    .A3(_07935_),
    .ZN(_08041_));
 OAI21_X1 _17312_ (.A(_07943_),
    .B1(_07916_),
    .B2(_07921_),
    .ZN(_08042_));
 AOI21_X1 _17313_ (.A(_06382_),
    .B1(_08041_),
    .B2(_08042_),
    .ZN(_08043_));
 AOI21_X2 _17314_ (.A(_07994_),
    .B1(_07910_),
    .B2(_07972_),
    .ZN(_08044_));
 AOI21_X1 _17315_ (.A(_08043_),
    .B1(_08044_),
    .B2(_08008_),
    .ZN(_08045_));
 NOR4_X4 _17316_ (.A1(_06338_),
    .A2(_06350_),
    .A3(_07914_),
    .A4(_07919_),
    .ZN(_08046_));
 NOR3_X2 _17317_ (.A1(_08007_),
    .A2(_07928_),
    .A3(_08046_),
    .ZN(_08047_));
 OR2_X1 _17318_ (.A1(_07994_),
    .A2(_08029_),
    .ZN(_08048_));
 AOI21_X1 _17319_ (.A(_08047_),
    .B1(_08048_),
    .B2(_08008_),
    .ZN(_08049_));
 BUF_X4 _17320_ (.A(_06425_),
    .Z(_08050_));
 MUX2_X1 _17321_ (.A(_08045_),
    .B(_08049_),
    .S(_08050_),
    .Z(_08051_));
 AOI211_X2 _17322_ (.A(_06447_),
    .B(_08040_),
    .C1(_08051_),
    .C2(_08034_),
    .ZN(_08052_));
 NOR3_X2 _17323_ (.A1(net1122),
    .A2(_07915_),
    .A3(_07920_),
    .ZN(_08053_));
 AOI221_X1 _17324_ (.A(_06350_),
    .B1(_06385_),
    .B2(_06397_),
    .C1(_07923_),
    .C2(_06401_),
    .ZN(_08054_));
 CLKBUF_X3 _17325_ (.A(_08054_),
    .Z(_08055_));
 OAI21_X1 _17326_ (.A(_07901_),
    .B1(_08053_),
    .B2(_08055_),
    .ZN(_08056_));
 BUF_X4 _17327_ (.A(_06425_),
    .Z(_08057_));
 AOI21_X1 _17328_ (.A(_08057_),
    .B1(_07928_),
    .B2(net39),
    .ZN(_08058_));
 NAND3_X2 _17329_ (.A1(_07913_),
    .A2(_07934_),
    .A3(_07935_),
    .ZN(_08059_));
 NAND3_X1 _17330_ (.A1(_07963_),
    .A2(_08059_),
    .A3(_07984_),
    .ZN(_08060_));
 OAI21_X1 _17331_ (.A(_08060_),
    .B1(_07999_),
    .B2(_07958_),
    .ZN(_08061_));
 AOI221_X2 _17332_ (.A(_06413_),
    .B1(_08056_),
    .B2(_08058_),
    .C1(_08061_),
    .C2(_08050_),
    .ZN(_08062_));
 AOI21_X1 _17333_ (.A(_07957_),
    .B1(_08059_),
    .B2(_07984_),
    .ZN(_08063_));
 XNOR2_X1 _17334_ (.A(net39),
    .B(_07911_),
    .ZN(_08064_));
 BUF_X4 _17335_ (.A(_07950_),
    .Z(_08065_));
 AOI211_X2 _17336_ (.A(_08050_),
    .B(_08063_),
    .C1(_08064_),
    .C2(_08065_),
    .ZN(_08066_));
 INV_X2 _17337_ (.A(_14735_),
    .ZN(_08067_));
 MUX2_X1 _17338_ (.A(_08067_),
    .B(net29),
    .S(_08008_),
    .Z(_08068_));
 CLKBUF_X3 _17339_ (.A(_07975_),
    .Z(_08069_));
 MUX2_X1 _17340_ (.A(_14747_),
    .B(_08068_),
    .S(_08069_),
    .Z(_08070_));
 BUF_X4 _17341_ (.A(_08050_),
    .Z(_08071_));
 AOI21_X1 _17342_ (.A(_08066_),
    .B1(_08070_),
    .B2(_08071_),
    .ZN(_08072_));
 AOI21_X1 _17343_ (.A(_08062_),
    .B1(_08072_),
    .B2(_00401_),
    .ZN(_08073_));
 AOI21_X1 _17344_ (.A(_08052_),
    .B1(_08073_),
    .B2(_00404_),
    .ZN(_08074_));
 NAND2_X4 _17345_ (.A1(_07900_),
    .A2(_07910_),
    .ZN(_08075_));
 AOI21_X1 _17346_ (.A(_08046_),
    .B1(_08069_),
    .B2(_07972_),
    .ZN(_08076_));
 OAI221_X2 _17347_ (.A(_06427_),
    .B1(_08075_),
    .B2(_07997_),
    .C1(_08076_),
    .C2(_14746_),
    .ZN(_08077_));
 BUF_X4 _17348_ (.A(_08057_),
    .Z(_08078_));
 NOR3_X4 _17349_ (.A1(_07905_),
    .A2(_07915_),
    .A3(_07920_),
    .ZN(_08079_));
 AOI21_X2 _17350_ (.A(_14742_),
    .B1(_07934_),
    .B2(_07935_),
    .ZN(_08080_));
 OAI21_X1 _17351_ (.A(_07974_),
    .B1(_08079_),
    .B2(_08080_),
    .ZN(_08081_));
 NOR3_X4 _17352_ (.A1(_08067_),
    .A2(_07915_),
    .A3(_07920_),
    .ZN(_08082_));
 OAI21_X1 _17353_ (.A(_08065_),
    .B1(_07994_),
    .B2(_08082_),
    .ZN(_08083_));
 NAND3_X1 _17354_ (.A1(_08078_),
    .A2(_08081_),
    .A3(_08083_),
    .ZN(_08084_));
 NAND3_X1 _17355_ (.A1(_08034_),
    .A2(_08077_),
    .A3(_08084_),
    .ZN(_08085_));
 AOI21_X1 _17356_ (.A(_08079_),
    .B1(_08069_),
    .B2(net1163),
    .ZN(_08086_));
 OAI221_X1 _17357_ (.A(_06427_),
    .B1(_08075_),
    .B2(_07961_),
    .C1(_08086_),
    .C2(_08065_),
    .ZN(_08087_));
 NOR3_X1 _17358_ (.A1(_06336_),
    .A2(net28),
    .A3(_07966_),
    .ZN(_08088_));
 XNOR2_X2 _17359_ (.A(net1168),
    .B(_06399_),
    .ZN(_08089_));
 NOR2_X4 _17360_ (.A1(_06380_),
    .A2(_06399_),
    .ZN(_08090_));
 AOI221_X2 _17361_ (.A(_08088_),
    .B1(_08089_),
    .B2(_06336_),
    .C1(_07940_),
    .C2(_08090_),
    .ZN(_08091_));
 CLKBUF_X3 _17362_ (.A(_06426_),
    .Z(_08092_));
 CLKBUF_X3 _17363_ (.A(_08092_),
    .Z(_08093_));
 OAI21_X1 _17364_ (.A(_08087_),
    .B1(_08091_),
    .B2(_08093_),
    .ZN(_08094_));
 OAI21_X1 _17365_ (.A(_08085_),
    .B1(_08094_),
    .B2(_00401_),
    .ZN(_08095_));
 OAI21_X1 _17366_ (.A(_08012_),
    .B1(_07966_),
    .B2(_07913_),
    .ZN(_08096_));
 AOI22_X1 _17367_ (.A1(_14732_),
    .A2(_08090_),
    .B1(_08096_),
    .B2(_07973_),
    .ZN(_08097_));
 OAI21_X1 _17368_ (.A(_07957_),
    .B1(_08046_),
    .B2(_08080_),
    .ZN(_08098_));
 OAI21_X1 _17369_ (.A(_08098_),
    .B1(_08048_),
    .B2(_07901_),
    .ZN(_08099_));
 MUX2_X1 _17370_ (.A(_08097_),
    .B(_08099_),
    .S(_08092_),
    .Z(_08100_));
 AOI21_X4 _17371_ (.A(net1118),
    .B1(_06385_),
    .B2(_06397_),
    .ZN(_08101_));
 OR3_X2 _17372_ (.A1(_07978_),
    .A2(_07900_),
    .A3(_08101_),
    .ZN(_08102_));
 NAND3_X1 _17373_ (.A1(_07961_),
    .A2(_07934_),
    .A3(_07935_),
    .ZN(_08103_));
 OAI21_X1 _17374_ (.A(_08103_),
    .B1(_07910_),
    .B2(_07968_),
    .ZN(_08104_));
 OAI21_X1 _17375_ (.A(_08102_),
    .B1(_08104_),
    .B2(_08008_),
    .ZN(_08105_));
 OAI21_X1 _17376_ (.A(_07957_),
    .B1(_07994_),
    .B2(_07978_),
    .ZN(_08106_));
 OAI21_X1 _17377_ (.A(_07936_),
    .B1(_06400_),
    .B2(_07968_),
    .ZN(_08107_));
 OAI21_X1 _17378_ (.A(_08106_),
    .B1(_08107_),
    .B2(_07901_),
    .ZN(_08108_));
 MUX2_X1 _17379_ (.A(_08105_),
    .B(_08108_),
    .S(_08092_),
    .Z(_08109_));
 MUX2_X1 _17380_ (.A(_08100_),
    .B(_08109_),
    .S(_06414_),
    .Z(_08110_));
 INV_X2 _17381_ (.A(_06447_),
    .ZN(_08111_));
 MUX2_X1 _17382_ (.A(_08095_),
    .B(_08110_),
    .S(_08111_),
    .Z(_08112_));
 MUX2_X1 _17383_ (.A(_08074_),
    .B(_08112_),
    .S(_00403_),
    .Z(_00017_));
 NOR2_X4 _17384_ (.A1(_06381_),
    .A2(_07907_),
    .ZN(_08113_));
 OR2_X1 _17385_ (.A1(_07978_),
    .A2(_08080_),
    .ZN(_08114_));
 AOI221_X1 _17386_ (.A(_08057_),
    .B1(_08113_),
    .B2(net1163),
    .C1(_08114_),
    .C2(_07974_),
    .ZN(_08115_));
 NAND3_X2 _17387_ (.A1(net1123),
    .A2(_07950_),
    .A3(_07975_),
    .ZN(_08116_));
 NAND2_X1 _17388_ (.A1(_14752_),
    .A2(_06400_),
    .ZN(_08117_));
 AOI21_X1 _17389_ (.A(_08093_),
    .B1(_08116_),
    .B2(_08117_),
    .ZN(_08118_));
 OAI21_X1 _17390_ (.A(_07948_),
    .B1(_08115_),
    .B2(_08118_),
    .ZN(_08119_));
 MUX2_X1 _17391_ (.A(_08003_),
    .B(_06352_),
    .S(_06382_),
    .Z(_08120_));
 MUX2_X1 _17392_ (.A(_14749_),
    .B(_08120_),
    .S(_00400_),
    .Z(_08121_));
 NAND3_X1 _17393_ (.A1(_06336_),
    .A2(_08007_),
    .A3(_07910_),
    .ZN(_08122_));
 OAI221_X1 _17394_ (.A(_08122_),
    .B1(_07944_),
    .B2(net99),
    .C1(_07961_),
    .C2(_07942_),
    .ZN(_08123_));
 MUX2_X1 _17395_ (.A(_08121_),
    .B(_08123_),
    .S(_08093_),
    .Z(_08124_));
 OAI21_X1 _17396_ (.A(_08119_),
    .B1(_08124_),
    .B2(_07948_),
    .ZN(_08125_));
 CLKBUF_X3 _17397_ (.A(_07973_),
    .Z(_08126_));
 AOI21_X1 _17398_ (.A(_08126_),
    .B1(_07933_),
    .B2(_08103_),
    .ZN(_08127_));
 NOR2_X1 _17399_ (.A1(net1119),
    .A2(_08002_),
    .ZN(_08128_));
 NOR4_X1 _17400_ (.A1(_08034_),
    .A2(_08071_),
    .A3(_08127_),
    .A4(_08128_),
    .ZN(_08129_));
 AOI21_X2 _17401_ (.A(_07983_),
    .B1(_07934_),
    .B2(_07935_),
    .ZN(_08130_));
 NOR3_X1 _17402_ (.A1(_08065_),
    .A2(_08046_),
    .A3(_08130_),
    .ZN(_08131_));
 NOR3_X1 _17403_ (.A1(_08126_),
    .A2(net1167),
    .A3(_08101_),
    .ZN(_08132_));
 NOR3_X1 _17404_ (.A1(_08093_),
    .A2(_08131_),
    .A3(_08132_),
    .ZN(_08133_));
 NOR3_X1 _17405_ (.A1(_07968_),
    .A2(_07916_),
    .A3(_07921_),
    .ZN(_08134_));
 NOR3_X1 _17406_ (.A1(_08126_),
    .A2(_08055_),
    .A3(_08134_),
    .ZN(_08135_));
 AND2_X1 _17407_ (.A1(_07955_),
    .A2(_08010_),
    .ZN(_08136_));
 AOI21_X1 _17408_ (.A(_08135_),
    .B1(_08136_),
    .B2(_14751_),
    .ZN(_08137_));
 AOI21_X1 _17409_ (.A(_08133_),
    .B1(_08137_),
    .B2(_00402_),
    .ZN(_08138_));
 AOI21_X1 _17410_ (.A(_08129_),
    .B1(_08138_),
    .B2(_00401_),
    .ZN(_08139_));
 NAND2_X1 _17411_ (.A1(_07904_),
    .A2(_08078_),
    .ZN(_08140_));
 MUX2_X1 _17412_ (.A(_08067_),
    .B(net1122),
    .S(_07974_),
    .Z(_08141_));
 AOI21_X1 _17413_ (.A(_08140_),
    .B1(_08141_),
    .B2(_00400_),
    .ZN(_08142_));
 NOR2_X1 _17414_ (.A1(net27),
    .A2(_07958_),
    .ZN(_08143_));
 NOR2_X1 _17415_ (.A1(_07913_),
    .A2(_06382_),
    .ZN(_08144_));
 OAI21_X1 _17416_ (.A(_08069_),
    .B1(_08143_),
    .B2(_08144_),
    .ZN(_08145_));
 AOI21_X1 _17417_ (.A(_06448_),
    .B1(_08142_),
    .B2(_08145_),
    .ZN(_08146_));
 AOI22_X1 _17418_ (.A1(_00404_),
    .A2(_08125_),
    .B1(_08139_),
    .B2(_08146_),
    .ZN(_08147_));
 AOI21_X4 _17419_ (.A(_14740_),
    .B1(_06385_),
    .B2(_06397_),
    .ZN(_08148_));
 NOR2_X1 _17420_ (.A1(_07978_),
    .A2(_08148_),
    .ZN(_08149_));
 MUX2_X1 _17421_ (.A(_07995_),
    .B(_08149_),
    .S(_07963_),
    .Z(_08150_));
 AOI21_X1 _17422_ (.A(_08148_),
    .B1(_07910_),
    .B2(_06352_),
    .ZN(_08151_));
 MUX2_X1 _17423_ (.A(_07983_),
    .B(_08151_),
    .S(_06382_),
    .Z(_08152_));
 MUX2_X1 _17424_ (.A(_08150_),
    .B(_08152_),
    .S(_08057_),
    .Z(_08153_));
 NOR3_X1 _17425_ (.A1(_06381_),
    .A2(_08046_),
    .A3(_08101_),
    .ZN(_08154_));
 MUX2_X1 _17426_ (.A(_14740_),
    .B(net605),
    .S(_07907_),
    .Z(_08155_));
 AOI211_X2 _17427_ (.A(_06425_),
    .B(_08154_),
    .C1(_08155_),
    .C2(_06382_),
    .ZN(_08156_));
 NOR3_X1 _17428_ (.A1(_08008_),
    .A2(_08029_),
    .A3(_08101_),
    .ZN(_08157_));
 AOI21_X1 _17429_ (.A(_08148_),
    .B1(_07911_),
    .B2(_14732_),
    .ZN(_08158_));
 AOI21_X1 _17430_ (.A(_08157_),
    .B1(_08158_),
    .B2(_07974_),
    .ZN(_08159_));
 AOI21_X1 _17431_ (.A(_08156_),
    .B1(_08159_),
    .B2(_08078_),
    .ZN(_08160_));
 MUX2_X1 _17432_ (.A(_08153_),
    .B(_08160_),
    .S(_06414_),
    .Z(_08161_));
 NAND2_X1 _17433_ (.A1(_14754_),
    .A2(_07966_),
    .ZN(_08162_));
 NAND2_X1 _17434_ (.A1(_08007_),
    .A2(_08053_),
    .ZN(_08163_));
 NAND3_X1 _17435_ (.A1(_07903_),
    .A2(_08162_),
    .A3(_08163_),
    .ZN(_08164_));
 AOI21_X1 _17436_ (.A(_06411_),
    .B1(_07910_),
    .B2(_14749_),
    .ZN(_08165_));
 NAND2_X1 _17437_ (.A1(_08022_),
    .A2(_08165_),
    .ZN(_08166_));
 AOI21_X4 _17438_ (.A(_07913_),
    .B1(_07934_),
    .B2(_07935_),
    .ZN(_08167_));
 OAI21_X1 _17439_ (.A(_08167_),
    .B1(_06412_),
    .B2(_14754_),
    .ZN(_08168_));
 OAI21_X1 _17440_ (.A(_07978_),
    .B1(_06411_),
    .B2(_14749_),
    .ZN(_08169_));
 NAND2_X1 _17441_ (.A1(_08168_),
    .A2(_08169_),
    .ZN(_08170_));
 AOI221_X2 _17442_ (.A(_08057_),
    .B1(_08164_),
    .B2(_08166_),
    .C1(_08170_),
    .C2(_07958_),
    .ZN(_08171_));
 MUX2_X1 _17443_ (.A(_06336_),
    .B(_08007_),
    .S(net28),
    .Z(_08172_));
 MUX2_X1 _17444_ (.A(_14756_),
    .B(_08172_),
    .S(_07911_),
    .Z(_08173_));
 OAI22_X2 _17445_ (.A1(_06338_),
    .A2(_06350_),
    .B1(_07916_),
    .B2(_07921_),
    .ZN(_08174_));
 AND3_X1 _17446_ (.A1(_07973_),
    .A2(_08174_),
    .A3(_08009_),
    .ZN(_08175_));
 AOI21_X1 _17447_ (.A(_08175_),
    .B1(_08114_),
    .B2(_07958_),
    .ZN(_08176_));
 MUX2_X1 _17448_ (.A(_08173_),
    .B(_08176_),
    .S(_06413_),
    .Z(_08177_));
 AOI21_X1 _17449_ (.A(_08171_),
    .B1(_08177_),
    .B2(_08071_),
    .ZN(_08178_));
 MUX2_X1 _17450_ (.A(_08161_),
    .B(_08178_),
    .S(_00404_),
    .Z(_08179_));
 MUX2_X1 _17451_ (.A(_08147_),
    .B(_08179_),
    .S(_00403_),
    .Z(_00018_));
 NOR3_X1 _17452_ (.A1(_07943_),
    .A2(_07916_),
    .A3(_07921_),
    .ZN(_08180_));
 AOI21_X4 _17453_ (.A(_14738_),
    .B1(_07934_),
    .B2(_07935_),
    .ZN(_08181_));
 NOR3_X1 _17454_ (.A1(_14746_),
    .A2(_08180_),
    .A3(_08181_),
    .ZN(_08182_));
 NOR3_X1 _17455_ (.A1(_14751_),
    .A2(_07994_),
    .A3(_08079_),
    .ZN(_08183_));
 NOR3_X1 _17456_ (.A1(_08071_),
    .A2(_08182_),
    .A3(_08183_),
    .ZN(_08184_));
 OR2_X1 _17457_ (.A1(_14749_),
    .A2(_07911_),
    .ZN(_08185_));
 NOR2_X1 _17458_ (.A1(_06336_),
    .A2(_07957_),
    .ZN(_08186_));
 OAI22_X1 _17459_ (.A1(_07940_),
    .A2(_08075_),
    .B1(_08185_),
    .B2(_08186_),
    .ZN(_08187_));
 OAI21_X1 _17460_ (.A(_08034_),
    .B1(_00402_),
    .B2(_08187_),
    .ZN(_08188_));
 NOR2_X1 _17461_ (.A1(_07994_),
    .A2(_08046_),
    .ZN(_08189_));
 OAI221_X1 _17462_ (.A(_07941_),
    .B1(_08189_),
    .B2(_08126_),
    .C1(_08174_),
    .C2(_07902_),
    .ZN(_08190_));
 NOR3_X1 _17463_ (.A1(_08065_),
    .A2(_07998_),
    .A3(_08167_),
    .ZN(_08191_));
 NOR3_X1 _17464_ (.A1(_07974_),
    .A2(_08082_),
    .A3(_08055_),
    .ZN(_08192_));
 NOR2_X1 _17465_ (.A1(_08191_),
    .A2(_08192_),
    .ZN(_08193_));
 MUX2_X1 _17466_ (.A(_08190_),
    .B(_08193_),
    .S(_08093_),
    .Z(_08194_));
 OAI221_X1 _17467_ (.A(_00404_),
    .B1(_08184_),
    .B2(_08188_),
    .C1(_08194_),
    .C2(_00401_),
    .ZN(_08195_));
 NAND3_X1 _17468_ (.A1(net39),
    .A2(_07963_),
    .A3(_07966_),
    .ZN(_08196_));
 NAND4_X1 _17469_ (.A1(_07903_),
    .A2(_08057_),
    .A3(_08122_),
    .A4(_08196_),
    .ZN(_08197_));
 OAI21_X1 _17470_ (.A(_07955_),
    .B1(_07973_),
    .B2(_06336_),
    .ZN(_08198_));
 AOI21_X1 _17471_ (.A(_08021_),
    .B1(_07901_),
    .B2(_14732_),
    .ZN(_08199_));
 AOI221_X2 _17472_ (.A(_08197_),
    .B1(_08198_),
    .B2(net1121),
    .C1(_07940_),
    .C2(_08199_),
    .ZN(_08200_));
 OAI21_X1 _17473_ (.A(_07900_),
    .B1(_08079_),
    .B2(_08181_),
    .ZN(_08201_));
 OAI21_X1 _17474_ (.A(_08201_),
    .B1(_07908_),
    .B2(net28),
    .ZN(_08202_));
 INV_X1 _17475_ (.A(_07968_),
    .ZN(_08203_));
 OAI22_X1 _17476_ (.A1(_08203_),
    .A2(_07967_),
    .B1(_08057_),
    .B2(_08010_),
    .ZN(_08204_));
 AOI221_X1 _17477_ (.A(_07903_),
    .B1(_08057_),
    .B2(_08202_),
    .C1(_08204_),
    .C2(_07974_),
    .ZN(_08205_));
 NAND3_X1 _17478_ (.A1(net829),
    .A2(_06383_),
    .A3(_07967_),
    .ZN(_08206_));
 INV_X1 _17479_ (.A(_07981_),
    .ZN(_08207_));
 OAI21_X1 _17480_ (.A(_08206_),
    .B1(_08089_),
    .B2(_08207_),
    .ZN(_08208_));
 NOR3_X1 _17481_ (.A1(_08034_),
    .A2(_08078_),
    .A3(_08208_),
    .ZN(_08209_));
 OR3_X1 _17482_ (.A1(_08200_),
    .A2(_08205_),
    .A3(_08209_),
    .ZN(_08210_));
 OAI21_X1 _17483_ (.A(_08195_),
    .B1(_08210_),
    .B2(_00404_),
    .ZN(_08211_));
 NAND2_X1 _17484_ (.A1(_06351_),
    .A2(_06399_),
    .ZN(_08212_));
 NOR2_X2 _17485_ (.A1(_06411_),
    .A2(_06425_),
    .ZN(_08213_));
 AOI211_X2 _17486_ (.A(net1168),
    .B(_08212_),
    .C1(_08213_),
    .C2(net602),
    .ZN(_08214_));
 NOR2_X1 _17487_ (.A1(_06411_),
    .A2(_06426_),
    .ZN(_08215_));
 AOI21_X1 _17488_ (.A(_07998_),
    .B1(_07907_),
    .B2(_07981_),
    .ZN(_08216_));
 OAI21_X1 _17489_ (.A(_08215_),
    .B1(_08216_),
    .B2(_07973_),
    .ZN(_08217_));
 NOR2_X1 _17490_ (.A1(_08021_),
    .A2(_08181_),
    .ZN(_08218_));
 OAI221_X2 _17491_ (.A(_08213_),
    .B1(_08218_),
    .B2(_08007_),
    .C1(_08212_),
    .C2(net1209),
    .ZN(_08219_));
 AOI221_X2 _17492_ (.A(_08214_),
    .B1(_08217_),
    .B2(_08219_),
    .C1(_08167_),
    .C2(_07974_),
    .ZN(_08220_));
 MUX2_X1 _17493_ (.A(net28),
    .B(_08007_),
    .S(net603),
    .Z(_08221_));
 AOI221_X2 _17494_ (.A(_06426_),
    .B1(_08113_),
    .B2(net1122),
    .C1(_08221_),
    .C2(_07967_),
    .ZN(_08222_));
 NAND3_X1 _17495_ (.A1(_08126_),
    .A2(_08009_),
    .A3(_08012_),
    .ZN(_08223_));
 AOI21_X1 _17496_ (.A(_08053_),
    .B1(_08069_),
    .B2(_07940_),
    .ZN(_08224_));
 OAI21_X1 _17497_ (.A(_08223_),
    .B1(_08224_),
    .B2(_14751_),
    .ZN(_08225_));
 AOI21_X1 _17498_ (.A(_08222_),
    .B1(_08225_),
    .B2(_08093_),
    .ZN(_08226_));
 AOI21_X1 _17499_ (.A(_08220_),
    .B1(_08226_),
    .B2(_07948_),
    .ZN(_08227_));
 OAI21_X1 _17500_ (.A(_07955_),
    .B1(_06399_),
    .B2(_07960_),
    .ZN(_08228_));
 NAND3_X4 _17501_ (.A1(_14740_),
    .A2(_06385_),
    .A3(_06397_),
    .ZN(_08229_));
 OAI21_X4 _17502_ (.A(_08229_),
    .B1(_06399_),
    .B2(_14738_),
    .ZN(_08230_));
 MUX2_X1 _17503_ (.A(_08228_),
    .B(_08230_),
    .S(_07963_),
    .Z(_08231_));
 OAI21_X1 _17504_ (.A(net39),
    .B1(_07963_),
    .B2(_07928_),
    .ZN(_08232_));
 OAI221_X1 _17505_ (.A(_08232_),
    .B1(_07944_),
    .B2(net98),
    .C1(_07943_),
    .C2(_08002_),
    .ZN(_08233_));
 MUX2_X1 _17506_ (.A(_08231_),
    .B(_08233_),
    .S(_08092_),
    .Z(_08234_));
 AOI21_X1 _17507_ (.A(_08101_),
    .B1(_08021_),
    .B2(_08092_),
    .ZN(_08235_));
 NAND2_X1 _17508_ (.A1(_06336_),
    .A2(_07907_),
    .ZN(_08236_));
 NAND2_X1 _17509_ (.A1(_08229_),
    .A2(_08023_),
    .ZN(_08237_));
 MUX2_X1 _17510_ (.A(_08236_),
    .B(_08237_),
    .S(_06426_),
    .Z(_08238_));
 MUX2_X1 _17511_ (.A(_08235_),
    .B(_08238_),
    .S(_06383_),
    .Z(_08239_));
 MUX2_X1 _17512_ (.A(_08234_),
    .B(_08239_),
    .S(_06414_),
    .Z(_08240_));
 MUX2_X1 _17513_ (.A(_08227_),
    .B(_08240_),
    .S(_08111_),
    .Z(_08241_));
 MUX2_X2 _17514_ (.A(_08211_),
    .B(_08241_),
    .S(_00403_),
    .Z(_00019_));
 AOI21_X1 _17515_ (.A(_08046_),
    .B1(_07907_),
    .B2(_07983_),
    .ZN(_08242_));
 OAI21_X1 _17516_ (.A(_07937_),
    .B1(_08242_),
    .B2(_06382_),
    .ZN(_08243_));
 NOR2_X1 _17517_ (.A1(_08004_),
    .A2(_08101_),
    .ZN(_08244_));
 MUX2_X1 _17518_ (.A(_08244_),
    .B(_08237_),
    .S(_07900_),
    .Z(_08245_));
 MUX2_X1 _17519_ (.A(_08243_),
    .B(_08245_),
    .S(_08092_),
    .Z(_08246_));
 NAND2_X1 _17520_ (.A1(_08207_),
    .A2(_06382_),
    .ZN(_08247_));
 AOI21_X1 _17521_ (.A(_06425_),
    .B1(_08060_),
    .B2(_08247_),
    .ZN(_08248_));
 NOR3_X1 _17522_ (.A1(_07963_),
    .A2(net1166),
    .A3(_08130_),
    .ZN(_08249_));
 AOI21_X1 _17523_ (.A(_08101_),
    .B1(_06400_),
    .B2(_06352_),
    .ZN(_08250_));
 AOI21_X1 _17524_ (.A(_08249_),
    .B1(_08250_),
    .B2(_07901_),
    .ZN(_08251_));
 AOI21_X1 _17525_ (.A(_08248_),
    .B1(_08251_),
    .B2(_08050_),
    .ZN(_08252_));
 MUX2_X1 _17526_ (.A(_08246_),
    .B(_08252_),
    .S(_06413_),
    .Z(_08253_));
 NAND2_X2 _17527_ (.A1(_06352_),
    .A2(_06381_),
    .ZN(_08254_));
 OAI21_X1 _17528_ (.A(_07966_),
    .B1(_06412_),
    .B2(_07968_),
    .ZN(_08255_));
 OAI21_X1 _17529_ (.A(_08057_),
    .B1(_08254_),
    .B2(_08255_),
    .ZN(_08256_));
 MUX2_X1 _17530_ (.A(_07981_),
    .B(_06336_),
    .S(_08007_),
    .Z(_08257_));
 NOR2_X2 _17531_ (.A1(_07966_),
    .A2(_06411_),
    .ZN(_08258_));
 MUX2_X1 _17532_ (.A(_08203_),
    .B(_07943_),
    .S(net1168),
    .Z(_08259_));
 OAI22_X2 _17533_ (.A1(net27),
    .A2(_07955_),
    .B1(_08259_),
    .B2(_07911_),
    .ZN(_08260_));
 AOI221_X2 _17534_ (.A(_08256_),
    .B1(_08257_),
    .B2(_08258_),
    .C1(_07903_),
    .C2(_08260_),
    .ZN(_08261_));
 AOI22_X1 _17535_ (.A1(_00400_),
    .A2(_07903_),
    .B1(_08055_),
    .B2(_07968_),
    .ZN(_08262_));
 NOR2_X1 _17536_ (.A1(_14746_),
    .A2(_08262_),
    .ZN(_08263_));
 OAI21_X1 _17537_ (.A(_07904_),
    .B1(_14751_),
    .B2(_07943_),
    .ZN(_08264_));
 AOI21_X1 _17538_ (.A(_08263_),
    .B1(_08264_),
    .B2(_08055_),
    .ZN(_08265_));
 OAI21_X1 _17539_ (.A(_08261_),
    .B1(_08265_),
    .B2(_14732_),
    .ZN(_08266_));
 OAI21_X1 _17540_ (.A(_06383_),
    .B1(_07996_),
    .B2(_08046_),
    .ZN(_08267_));
 AOI21_X1 _17541_ (.A(_07904_),
    .B1(_08017_),
    .B2(_08267_),
    .ZN(_08268_));
 AOI221_X1 _17542_ (.A(_06412_),
    .B1(_08113_),
    .B2(_07913_),
    .C1(_07961_),
    .C2(_07975_),
    .ZN(_08269_));
 NOR3_X1 _17543_ (.A1(_08071_),
    .A2(_08268_),
    .A3(_08269_),
    .ZN(_08270_));
 NOR2_X1 _17544_ (.A1(_06448_),
    .A2(_08270_),
    .ZN(_08271_));
 AOI221_X2 _17545_ (.A(_06438_),
    .B1(_08253_),
    .B2(_06448_),
    .C1(_08266_),
    .C2(_08271_),
    .ZN(_08272_));
 NOR3_X1 _17546_ (.A1(_07958_),
    .A2(_08082_),
    .A3(_08080_),
    .ZN(_08273_));
 OAI21_X1 _17547_ (.A(_06414_),
    .B1(_08047_),
    .B2(_08273_),
    .ZN(_08274_));
 OAI22_X1 _17548_ (.A1(net49),
    .A2(_07908_),
    .B1(_08101_),
    .B2(_08126_),
    .ZN(_08275_));
 OAI21_X1 _17549_ (.A(_08274_),
    .B1(_08275_),
    .B2(_08034_),
    .ZN(_08276_));
 AOI21_X1 _17550_ (.A(_06413_),
    .B1(_07955_),
    .B2(net98),
    .ZN(_08277_));
 OAI221_X1 _17551_ (.A(_08277_),
    .B1(_08075_),
    .B2(_14737_),
    .C1(net49),
    .C2(_07908_),
    .ZN(_08278_));
 NOR2_X1 _17552_ (.A1(_08126_),
    .A2(_07936_),
    .ZN(_08279_));
 OAI21_X1 _17553_ (.A(_06414_),
    .B1(_08143_),
    .B2(_08279_),
    .ZN(_08280_));
 OAI21_X1 _17554_ (.A(_07994_),
    .B1(_14751_),
    .B2(net27),
    .ZN(_08281_));
 NAND3_X1 _17555_ (.A1(_08278_),
    .A2(_08280_),
    .A3(_08281_),
    .ZN(_08282_));
 MUX2_X1 _17556_ (.A(_08276_),
    .B(_08282_),
    .S(_06448_),
    .Z(_08283_));
 NOR2_X1 _17557_ (.A1(_08067_),
    .A2(_07957_),
    .ZN(_08284_));
 OAI21_X1 _17558_ (.A(_07967_),
    .B1(_08144_),
    .B2(_08284_),
    .ZN(_08285_));
 NOR2_X1 _17559_ (.A1(_07974_),
    .A2(_07903_),
    .ZN(_08286_));
 AOI221_X2 _17560_ (.A(_06447_),
    .B1(_07965_),
    .B2(_08285_),
    .C1(_08286_),
    .C2(_08104_),
    .ZN(_08287_));
 NAND2_X1 _17561_ (.A1(_14758_),
    .A2(_00400_),
    .ZN(_08288_));
 OAI221_X1 _17562_ (.A(_08288_),
    .B1(_08065_),
    .B2(_14732_),
    .C1(_07943_),
    .C2(_07944_),
    .ZN(_08289_));
 AOI21_X1 _17563_ (.A(_08018_),
    .B1(_08229_),
    .B2(_14746_),
    .ZN(_08290_));
 MUX2_X1 _17564_ (.A(_08289_),
    .B(_08290_),
    .S(_06414_),
    .Z(_08291_));
 AOI21_X1 _17565_ (.A(_08287_),
    .B1(_08291_),
    .B2(_00404_),
    .ZN(_08292_));
 MUX2_X1 _17566_ (.A(_08283_),
    .B(_08292_),
    .S(_00402_),
    .Z(_08293_));
 AOI21_X2 _17567_ (.A(_08272_),
    .B1(_08293_),
    .B2(_00403_),
    .ZN(_00020_));
 AOI222_X2 _17568_ (.A1(net829),
    .A2(_07928_),
    .B1(_08044_),
    .B2(_08008_),
    .C1(_08113_),
    .C2(net99),
    .ZN(_08294_));
 OAI21_X1 _17569_ (.A(_07968_),
    .B1(_07916_),
    .B2(_07921_),
    .ZN(_08295_));
 AOI21_X1 _17570_ (.A(_08126_),
    .B1(_08059_),
    .B2(_08295_),
    .ZN(_08296_));
 OAI21_X1 _17571_ (.A(_08050_),
    .B1(_07908_),
    .B2(net27),
    .ZN(_08297_));
 OAI221_X1 _17572_ (.A(_08034_),
    .B1(_08078_),
    .B2(_08294_),
    .C1(_08296_),
    .C2(_08297_),
    .ZN(_08298_));
 AOI21_X1 _17573_ (.A(_08180_),
    .B1(_08069_),
    .B2(net1120),
    .ZN(_08299_));
 OAI221_X1 _17574_ (.A(_08050_),
    .B1(_08002_),
    .B2(_07940_),
    .C1(_08299_),
    .C2(_14751_),
    .ZN(_08300_));
 AOI22_X1 _17575_ (.A1(net98),
    .A2(_07944_),
    .B1(_08055_),
    .B2(net829),
    .ZN(_08301_));
 OAI21_X1 _17576_ (.A(_08300_),
    .B1(_08301_),
    .B2(_08071_),
    .ZN(_08302_));
 OAI21_X1 _17577_ (.A(_08298_),
    .B1(_08302_),
    .B2(_00401_),
    .ZN(_08303_));
 NOR2_X1 _17578_ (.A1(_08065_),
    .A2(_08228_),
    .ZN(_08304_));
 NAND2_X1 _17579_ (.A1(_06427_),
    .A2(_08116_),
    .ZN(_08305_));
 OAI21_X1 _17580_ (.A(_08009_),
    .B1(_07962_),
    .B2(_00400_),
    .ZN(_08306_));
 OAI22_X1 _17581_ (.A1(_08304_),
    .A2(_08305_),
    .B1(_08306_),
    .B2(_06427_),
    .ZN(_08307_));
 NAND2_X1 _17582_ (.A1(_07997_),
    .A2(_07900_),
    .ZN(_08308_));
 AOI221_X2 _17583_ (.A(_06425_),
    .B1(_08090_),
    .B2(_07983_),
    .C1(_08308_),
    .C2(_07910_),
    .ZN(_08309_));
 AOI21_X1 _17584_ (.A(_07950_),
    .B1(_08059_),
    .B2(_08010_),
    .ZN(_08310_));
 OAI21_X1 _17585_ (.A(net1170),
    .B1(_07916_),
    .B2(_07921_),
    .ZN(_08311_));
 OAI21_X1 _17586_ (.A(_08311_),
    .B1(_07975_),
    .B2(_14738_),
    .ZN(_08312_));
 AOI21_X1 _17587_ (.A(_08310_),
    .B1(_08312_),
    .B2(_07958_),
    .ZN(_08313_));
 AOI21_X1 _17588_ (.A(_08309_),
    .B1(_08313_),
    .B2(_08078_),
    .ZN(_08314_));
 MUX2_X1 _17589_ (.A(_08307_),
    .B(_08314_),
    .S(_06414_),
    .Z(_08315_));
 MUX2_X1 _17590_ (.A(_08303_),
    .B(_08315_),
    .S(_08111_),
    .Z(_08316_));
 OAI21_X1 _17591_ (.A(_07950_),
    .B1(_07952_),
    .B2(_08055_),
    .ZN(_08317_));
 NAND3_X1 _17592_ (.A1(_08092_),
    .A2(_08030_),
    .A3(_08317_),
    .ZN(_08318_));
 NAND3_X1 _17593_ (.A1(_07973_),
    .A2(_08023_),
    .A3(_08229_),
    .ZN(_08319_));
 NAND2_X1 _17594_ (.A1(_07901_),
    .A2(_08021_),
    .ZN(_08320_));
 NAND3_X1 _17595_ (.A1(_08050_),
    .A2(_08319_),
    .A3(_08320_),
    .ZN(_08321_));
 AOI21_X1 _17596_ (.A(_06413_),
    .B1(_08318_),
    .B2(_08321_),
    .ZN(_08322_));
 AOI211_X2 _17597_ (.A(net1168),
    .B(_07996_),
    .C1(_06399_),
    .C2(_06336_),
    .ZN(_08323_));
 AOI21_X1 _17598_ (.A(_08082_),
    .B1(_07975_),
    .B2(_07981_),
    .ZN(_08324_));
 AOI21_X1 _17599_ (.A(_08323_),
    .B1(_08324_),
    .B2(_07901_),
    .ZN(_08325_));
 OAI21_X1 _17600_ (.A(_07984_),
    .B1(net1166),
    .B2(_08008_),
    .ZN(_08326_));
 MUX2_X1 _17601_ (.A(_08325_),
    .B(_08326_),
    .S(_08050_),
    .Z(_08327_));
 AOI211_X2 _17602_ (.A(_08111_),
    .B(_08322_),
    .C1(_08327_),
    .C2(_08034_),
    .ZN(_08328_));
 AOI21_X1 _17603_ (.A(_06400_),
    .B1(_07973_),
    .B2(_06336_),
    .ZN(_08329_));
 OAI21_X1 _17604_ (.A(_08329_),
    .B1(_06383_),
    .B2(net1163),
    .ZN(_08330_));
 AOI22_X2 _17605_ (.A1(_07972_),
    .A2(_07979_),
    .B1(_08312_),
    .B2(_07958_),
    .ZN(_08331_));
 AOI221_X2 _17606_ (.A(_06427_),
    .B1(_07965_),
    .B2(_08330_),
    .C1(_08331_),
    .C2(_06414_),
    .ZN(_08332_));
 NOR3_X1 _17607_ (.A1(_08065_),
    .A2(_07928_),
    .A3(_08079_),
    .ZN(_08333_));
 NOR3_X1 _17608_ (.A1(_08126_),
    .A2(net1167),
    .A3(_08148_),
    .ZN(_08334_));
 NOR3_X1 _17609_ (.A1(_07904_),
    .A2(_08333_),
    .A3(_08334_),
    .ZN(_08335_));
 OAI21_X1 _17610_ (.A(_08206_),
    .B1(_08055_),
    .B2(net49),
    .ZN(_08336_));
 AOI21_X1 _17611_ (.A(_08335_),
    .B1(_08336_),
    .B2(_07948_),
    .ZN(_08337_));
 AOI21_X1 _17612_ (.A(_08332_),
    .B1(_08337_),
    .B2(_00402_),
    .ZN(_08338_));
 AOI21_X1 _17613_ (.A(_08328_),
    .B1(_08338_),
    .B2(_08111_),
    .ZN(_08339_));
 MUX2_X2 _17614_ (.A(_08316_),
    .B(_08339_),
    .S(_00403_),
    .Z(_00021_));
 NOR2_X1 _17615_ (.A1(_06438_),
    .A2(_06447_),
    .ZN(_08340_));
 OAI221_X2 _17616_ (.A(_08215_),
    .B1(_08230_),
    .B2(_14751_),
    .C1(_08002_),
    .C2(net27),
    .ZN(_08341_));
 NAND2_X1 _17617_ (.A1(_08340_),
    .A2(_08341_),
    .ZN(_08342_));
 NAND3_X1 _17618_ (.A1(_07906_),
    .A2(_07973_),
    .A3(_07911_),
    .ZN(_08343_));
 OAI21_X1 _17619_ (.A(_07900_),
    .B1(_07994_),
    .B2(_07998_),
    .ZN(_08344_));
 AND2_X1 _17620_ (.A1(_06412_),
    .A2(_08344_),
    .ZN(_08345_));
 OAI21_X1 _17621_ (.A(_08254_),
    .B1(_08007_),
    .B2(_07981_),
    .ZN(_08346_));
 MUX2_X1 _17622_ (.A(_14748_),
    .B(_08346_),
    .S(_07966_),
    .Z(_08347_));
 AOI221_X2 _17623_ (.A(_08050_),
    .B1(_08345_),
    .B2(_08343_),
    .C1(_07903_),
    .C2(_08347_),
    .ZN(_08348_));
 OAI21_X1 _17624_ (.A(_08229_),
    .B1(_06400_),
    .B2(_07943_),
    .ZN(_08349_));
 AOI221_X2 _17625_ (.A(_06425_),
    .B1(_08113_),
    .B2(_07968_),
    .C1(_08349_),
    .C2(_08008_),
    .ZN(_08350_));
 NAND2_X1 _17626_ (.A1(_07940_),
    .A2(_08090_),
    .ZN(_08351_));
 OAI221_X1 _17627_ (.A(_08351_),
    .B1(_07942_),
    .B2(_14732_),
    .C1(_07981_),
    .C2(_08002_),
    .ZN(_08352_));
 AOI21_X1 _17628_ (.A(_08350_),
    .B1(_08352_),
    .B2(_08071_),
    .ZN(_08353_));
 NAND2_X1 _17629_ (.A1(_06438_),
    .A2(_06448_),
    .ZN(_08354_));
 OAI33_X1 _17630_ (.A1(_08142_),
    .A2(_08342_),
    .A3(_08348_),
    .B1(_08353_),
    .B2(_08354_),
    .B3(_07948_),
    .ZN(_08355_));
 MUX2_X1 _17631_ (.A(_07913_),
    .B(_08003_),
    .S(net1168),
    .Z(_08356_));
 OAI21_X1 _17632_ (.A(_08117_),
    .B1(_08356_),
    .B2(_07911_),
    .ZN(_08357_));
 NOR2_X1 _17633_ (.A1(net27),
    .A2(_07975_),
    .ZN(_08358_));
 OAI21_X1 _17634_ (.A(_07958_),
    .B1(_08358_),
    .B2(_08181_),
    .ZN(_08359_));
 AOI21_X1 _17635_ (.A(_08092_),
    .B1(_08053_),
    .B2(_06383_),
    .ZN(_08360_));
 AOI221_X2 _17636_ (.A(_07904_),
    .B1(_08092_),
    .B2(_08357_),
    .C1(_08359_),
    .C2(_08360_),
    .ZN(_08361_));
 NOR3_X1 _17637_ (.A1(_07901_),
    .A2(_08167_),
    .A3(_08046_),
    .ZN(_08362_));
 AOI21_X1 _17638_ (.A(_08362_),
    .B1(_08019_),
    .B2(_08065_),
    .ZN(_08363_));
 OAI221_X1 _17639_ (.A(_08163_),
    .B1(_07942_),
    .B2(net49),
    .C1(_07940_),
    .C2(_07944_),
    .ZN(_08364_));
 MUX2_X1 _17640_ (.A(_08363_),
    .B(_08364_),
    .S(_08078_),
    .Z(_08365_));
 AOI21_X1 _17641_ (.A(_08361_),
    .B1(_08365_),
    .B2(_07948_),
    .ZN(_08366_));
 NOR2_X1 _17642_ (.A1(_00403_),
    .A2(_08111_),
    .ZN(_08367_));
 AOI21_X1 _17643_ (.A(_07902_),
    .B1(net98),
    .B2(_06400_),
    .ZN(_08368_));
 OAI221_X1 _17644_ (.A(_06427_),
    .B1(_08186_),
    .B2(_08368_),
    .C1(_07908_),
    .C2(net1169),
    .ZN(_08369_));
 MUX2_X1 _17645_ (.A(net1122),
    .B(_06336_),
    .S(_06381_),
    .Z(_08370_));
 MUX2_X1 _17646_ (.A(_14747_),
    .B(_08370_),
    .S(_07967_),
    .Z(_08371_));
 OAI21_X1 _17647_ (.A(_08369_),
    .B1(_08371_),
    .B2(_06427_),
    .ZN(_08372_));
 AOI21_X1 _17648_ (.A(_08092_),
    .B1(_07955_),
    .B2(_07901_),
    .ZN(_08373_));
 NAND2_X1 _17649_ (.A1(_08319_),
    .A2(_08373_),
    .ZN(_08374_));
 AND2_X1 _17650_ (.A1(_07957_),
    .A2(_07955_),
    .ZN(_08375_));
 OAI221_X1 _17651_ (.A(_08116_),
    .B1(_08375_),
    .B2(net98),
    .C1(_08002_),
    .C2(_14732_),
    .ZN(_08376_));
 OAI21_X1 _17652_ (.A(_08374_),
    .B1(_08376_),
    .B2(_08078_),
    .ZN(_08377_));
 MUX2_X1 _17653_ (.A(_08372_),
    .B(_08377_),
    .S(_07904_),
    .Z(_08378_));
 AOI221_X2 _17654_ (.A(_08057_),
    .B1(_08075_),
    .B2(net98),
    .C1(_08046_),
    .C2(net49),
    .ZN(_08379_));
 NOR3_X1 _17655_ (.A1(_14746_),
    .A2(_08101_),
    .A3(_08134_),
    .ZN(_08380_));
 AOI21_X1 _17656_ (.A(_08148_),
    .B1(_00400_),
    .B2(_07961_),
    .ZN(_08381_));
 AOI21_X1 _17657_ (.A(_08380_),
    .B1(_08381_),
    .B2(_14746_),
    .ZN(_08382_));
 AOI21_X1 _17658_ (.A(_08379_),
    .B1(_08382_),
    .B2(_08071_),
    .ZN(_08383_));
 NAND2_X1 _17659_ (.A1(_07948_),
    .A2(_06448_),
    .ZN(_08384_));
 OAI22_X1 _17660_ (.A1(_00404_),
    .A2(_08378_),
    .B1(_08383_),
    .B2(_08384_),
    .ZN(_08385_));
 AOI221_X2 _17661_ (.A(_08355_),
    .B1(_08366_),
    .B2(_08367_),
    .C1(_08385_),
    .C2(_00403_),
    .ZN(_00022_));
 NAND3_X1 _17662_ (.A1(_06383_),
    .A2(_07967_),
    .A3(_07903_),
    .ZN(_08386_));
 AOI21_X1 _17663_ (.A(net98),
    .B1(_08075_),
    .B2(_08386_),
    .ZN(_08387_));
 NAND2_X1 _17664_ (.A1(_06400_),
    .A2(_06412_),
    .ZN(_08388_));
 OAI33_X1 _17665_ (.A1(_07961_),
    .A2(_06413_),
    .A3(_07944_),
    .B1(_08388_),
    .B2(_07950_),
    .B3(_07902_),
    .ZN(_08389_));
 NAND3_X1 _17666_ (.A1(_14737_),
    .A2(_07911_),
    .A3(_07903_),
    .ZN(_08390_));
 NAND2_X1 _17667_ (.A1(_07967_),
    .A2(_06413_),
    .ZN(_08391_));
 AOI21_X1 _17668_ (.A(_14732_),
    .B1(_08390_),
    .B2(_08391_),
    .ZN(_08392_));
 NOR4_X1 _17669_ (.A1(_08078_),
    .A2(_08387_),
    .A3(_08389_),
    .A4(_08392_),
    .ZN(_08393_));
 OAI21_X1 _17670_ (.A(_07961_),
    .B1(_08090_),
    .B2(_07976_),
    .ZN(_08394_));
 AOI221_X1 _17671_ (.A(_07950_),
    .B1(_07975_),
    .B2(_07913_),
    .C1(_08258_),
    .C2(net1122),
    .ZN(_08395_));
 OAI21_X1 _17672_ (.A(_08394_),
    .B1(_08395_),
    .B2(_08286_),
    .ZN(_08396_));
 AOI21_X1 _17673_ (.A(_08393_),
    .B1(_08396_),
    .B2(_08071_),
    .ZN(_08397_));
 NAND4_X1 _17674_ (.A1(_08078_),
    .A2(_08343_),
    .A3(_08106_),
    .A4(_08162_),
    .ZN(_08398_));
 NOR3_X1 _17675_ (.A1(_07958_),
    .A2(_07996_),
    .A3(_08082_),
    .ZN(_08399_));
 OAI21_X1 _17676_ (.A(_08093_),
    .B1(_08047_),
    .B2(_08399_),
    .ZN(_08400_));
 NAND3_X1 _17677_ (.A1(_08034_),
    .A2(_08398_),
    .A3(_08400_),
    .ZN(_08401_));
 OAI221_X1 _17678_ (.A(_06427_),
    .B1(_07944_),
    .B2(_08203_),
    .C1(_07961_),
    .C2(_08069_),
    .ZN(_08402_));
 MUX2_X1 _17679_ (.A(_07940_),
    .B(_08207_),
    .S(_08008_),
    .Z(_08403_));
 OAI21_X1 _17680_ (.A(_08288_),
    .B1(_08403_),
    .B2(_00400_),
    .ZN(_08404_));
 OAI21_X1 _17681_ (.A(_08402_),
    .B1(_08404_),
    .B2(_08093_),
    .ZN(_08405_));
 OAI21_X1 _17682_ (.A(_08401_),
    .B1(_08405_),
    .B2(_00401_),
    .ZN(_08406_));
 MUX2_X1 _17683_ (.A(_08397_),
    .B(_08406_),
    .S(_06448_),
    .Z(_08407_));
 NOR2_X1 _17684_ (.A1(_07943_),
    .A2(_08065_),
    .ZN(_08408_));
 OAI21_X1 _17685_ (.A(_08295_),
    .B1(_08069_),
    .B2(net27),
    .ZN(_08409_));
 AOI21_X1 _17686_ (.A(_08408_),
    .B1(_08409_),
    .B2(_14746_),
    .ZN(_08410_));
 NOR2_X1 _17687_ (.A1(_00402_),
    .A2(_08410_),
    .ZN(_08411_));
 NAND3_X1 _17688_ (.A1(_14746_),
    .A2(_08009_),
    .A3(_08012_),
    .ZN(_08412_));
 AOI21_X1 _17689_ (.A(_08071_),
    .B1(_08081_),
    .B2(_08412_),
    .ZN(_08413_));
 NOR3_X1 _17690_ (.A1(_00401_),
    .A2(_08411_),
    .A3(_08413_),
    .ZN(_08414_));
 AOI21_X1 _17691_ (.A(_08069_),
    .B1(net27),
    .B2(net49),
    .ZN(_08415_));
 AOI21_X1 _17692_ (.A(_08130_),
    .B1(_08254_),
    .B2(_08415_),
    .ZN(_08416_));
 NOR3_X1 _17693_ (.A1(_07948_),
    .A2(_00402_),
    .A3(_08416_),
    .ZN(_08417_));
 NAND2_X1 _17694_ (.A1(_00401_),
    .A2(_00402_),
    .ZN(_08418_));
 OAI21_X1 _17695_ (.A(_08254_),
    .B1(_08126_),
    .B2(_07961_),
    .ZN(_08419_));
 MUX2_X1 _17696_ (.A(_08257_),
    .B(_08419_),
    .S(_08069_),
    .Z(_08420_));
 OAI21_X1 _17697_ (.A(_06448_),
    .B1(_08418_),
    .B2(_08420_),
    .ZN(_08421_));
 OAI221_X1 _17698_ (.A(_06427_),
    .B1(_08075_),
    .B2(_07981_),
    .C1(_08250_),
    .C2(_14746_),
    .ZN(_08422_));
 AND2_X1 _17699_ (.A1(_14749_),
    .A2(_07910_),
    .ZN(_08423_));
 OAI21_X1 _17700_ (.A(_08311_),
    .B1(_07966_),
    .B2(_06336_),
    .ZN(_08424_));
 AOI221_X2 _17701_ (.A(_08423_),
    .B1(_08424_),
    .B2(_07973_),
    .C1(_08090_),
    .C2(_07981_),
    .ZN(_08425_));
 OAI21_X1 _17702_ (.A(_08422_),
    .B1(_08425_),
    .B2(_00402_),
    .ZN(_08426_));
 NOR2_X1 _17703_ (.A1(_00401_),
    .A2(_08426_),
    .ZN(_08427_));
 NOR2_X1 _17704_ (.A1(net829),
    .A2(_07944_),
    .ZN(_08428_));
 NOR2_X1 _17705_ (.A1(_07940_),
    .A2(_07942_),
    .ZN(_08429_));
 NOR4_X1 _17706_ (.A1(_08093_),
    .A2(_08428_),
    .A3(_08128_),
    .A4(_08429_),
    .ZN(_08430_));
 OAI21_X1 _17707_ (.A(_07937_),
    .B1(_08044_),
    .B2(_07974_),
    .ZN(_08431_));
 AND2_X1 _17708_ (.A1(_08093_),
    .A2(_08431_),
    .ZN(_08432_));
 NOR3_X1 _17709_ (.A1(_07948_),
    .A2(_08430_),
    .A3(_08432_),
    .ZN(_08433_));
 OAI33_X1 _17710_ (.A1(_08414_),
    .A2(_08417_),
    .A3(_08421_),
    .B1(_08427_),
    .B2(_08433_),
    .B3(_00404_),
    .ZN(_08434_));
 MUX2_X2 _17711_ (.A(_08407_),
    .B(_08434_),
    .S(_00403_),
    .Z(_00023_));
 BUF_X8 _17712_ (.A(_06626_),
    .Z(_08435_));
 BUF_X16 _17713_ (.A(_08435_),
    .Z(_14760_));
 CLKBUF_X3 _17714_ (.A(_06642_),
    .Z(_08436_));
 BUF_X4 _17715_ (.A(_08436_),
    .Z(_08437_));
 BUF_X4 _17716_ (.A(_08437_),
    .Z(_08438_));
 BUF_X4 _17717_ (.A(_08438_),
    .Z(_14780_));
 BUF_X8 _17718_ (.A(_06610_),
    .Z(_14761_));
 AND2_X2 _17719_ (.A1(net18),
    .A2(net81),
    .ZN(_08439_));
 NOR2_X1 _17720_ (.A1(net6),
    .A2(_06633_),
    .ZN(_08440_));
 NOR2_X1 _17721_ (.A1(net6),
    .A2(_06631_),
    .ZN(_08441_));
 MUX2_X2 _17722_ (.A(_08440_),
    .B(_08441_),
    .S(_06640_),
    .Z(_08442_));
 NOR4_X4 _17723_ (.A1(_08439_),
    .A2(_08442_),
    .A3(_06647_),
    .A4(_06661_),
    .ZN(_08443_));
 BUF_X2 clone51 (.A(net504),
    .Z(net51));
 INV_X1 _17725_ (.A(net1001),
    .ZN(_08445_));
 CLKBUF_X3 _17726_ (.A(_14778_),
    .Z(_08446_));
 BUF_X4 _17727_ (.A(_06648_),
    .Z(_08447_));
 BUF_X4 _17728_ (.A(_06661_),
    .Z(_08448_));
 BUF_X4 _17729_ (.A(_08448_),
    .Z(_08449_));
 OAI21_X2 _17730_ (.A(_08446_),
    .B1(_08447_),
    .B2(_08449_),
    .ZN(_08450_));
 BUF_X1 rebuffer664 (.A(_15093_),
    .Z(net1127));
 BUF_X8 _17732_ (.A(net791),
    .Z(_08452_));
 OAI21_X2 _17733_ (.A(_08450_),
    .B1(_06663_),
    .B2(_08452_),
    .ZN(_08453_));
 AOI221_X2 _17734_ (.A(_06692_),
    .B1(_08443_),
    .B2(_08445_),
    .C1(_08437_),
    .C2(_08453_),
    .ZN(_08454_));
 BUF_X4 _17735_ (.A(_14763_),
    .Z(_08455_));
 AND2_X1 _17736_ (.A1(_08455_),
    .A2(_08443_),
    .ZN(_08456_));
 AOI21_X1 _17737_ (.A(_08456_),
    .B1(_00395_),
    .B2(_14783_),
    .ZN(_08457_));
 BUF_X4 _17738_ (.A(_06692_),
    .Z(_08458_));
 CLKBUF_X3 _17739_ (.A(_08458_),
    .Z(_08459_));
 AOI21_X2 _17740_ (.A(_08454_),
    .B1(_08457_),
    .B2(_08459_),
    .ZN(_08460_));
 NAND2_X4 _17741_ (.A1(_06245_),
    .A2(_06646_),
    .ZN(_08461_));
 NAND2_X1 _17742_ (.A1(_06217_),
    .A2(_06652_),
    .ZN(_08462_));
 NAND2_X1 _17743_ (.A1(_06217_),
    .A2(_06650_),
    .ZN(_08463_));
 MUX2_X2 _17744_ (.A(_08462_),
    .B(_08463_),
    .S(_06659_),
    .Z(_08464_));
 BUF_X8 _17745_ (.A(_08464_),
    .Z(_08465_));
 AOI221_X2 _17746_ (.A(_08442_),
    .B1(_08461_),
    .B2(_08465_),
    .C1(net81),
    .C2(_06279_),
    .ZN(_08466_));
 BUF_X4 _17747_ (.A(_08466_),
    .Z(_08467_));
 BUF_X4 _17748_ (.A(_14774_),
    .Z(_08468_));
 INV_X4 _17749_ (.A(net1230),
    .ZN(_08469_));
 OAI21_X4 _17750_ (.A(_08469_),
    .B1(_06648_),
    .B2(_08448_),
    .ZN(_08470_));
 NAND3_X2 _17751_ (.A1(_08446_),
    .A2(_08461_),
    .A3(_08465_),
    .ZN(_08471_));
 NAND2_X1 _17752_ (.A1(_08470_),
    .A2(_08471_),
    .ZN(_08472_));
 AOI221_X2 _17753_ (.A(_06692_),
    .B1(_08467_),
    .B2(_08468_),
    .C1(_08472_),
    .C2(_08437_),
    .ZN(_08473_));
 BUF_X4 _17754_ (.A(_06643_),
    .Z(_08474_));
 NOR3_X1 _17755_ (.A1(net1230),
    .A2(_08447_),
    .A3(_08449_),
    .ZN(_08475_));
 NOR2_X4 clone100 (.A1(_05530_),
    .A2(net528),
    .ZN(net100));
 AOI21_X2 _17757_ (.A(net789),
    .B1(_08461_),
    .B2(_08465_),
    .ZN(_08477_));
 OR3_X2 _17758_ (.A1(_08477_),
    .A2(_08475_),
    .A3(_08474_),
    .ZN(_08478_));
 BUF_X4 _17759_ (.A(_06662_),
    .Z(_08479_));
 BUF_X4 _17760_ (.A(_08479_),
    .Z(_08480_));
 XNOR2_X1 _17761_ (.A(net1116),
    .B(_08480_),
    .ZN(_08481_));
 BUF_X4 _17762_ (.A(_08436_),
    .Z(_08482_));
 BUF_X4 _17763_ (.A(_08482_),
    .Z(_08483_));
 OAI21_X1 _17764_ (.A(_08478_),
    .B1(_08481_),
    .B2(_08483_),
    .ZN(_08484_));
 AOI21_X1 _17765_ (.A(_08473_),
    .B1(_08484_),
    .B2(_08459_),
    .ZN(_08485_));
 BUF_X4 _17766_ (.A(_06677_),
    .Z(_08486_));
 CLKBUF_X3 _17767_ (.A(_08486_),
    .Z(_08487_));
 MUX2_X1 _17768_ (.A(_08460_),
    .B(_08485_),
    .S(_08487_),
    .Z(_08488_));
 AOI21_X4 _17769_ (.A(net1001),
    .B1(_08461_),
    .B2(_08465_),
    .ZN(_08489_));
 BUF_X8 _17770_ (.A(_08455_),
    .Z(_08490_));
 AOI221_X2 _17771_ (.A(_08489_),
    .B1(_06641_),
    .B2(_06629_),
    .C1(_08490_),
    .C2(_06662_),
    .ZN(_08491_));
 BUF_X2 _17772_ (.A(_14762_),
    .Z(_08492_));
 NOR3_X4 _17773_ (.A1(_08492_),
    .A2(_06648_),
    .A3(_08448_),
    .ZN(_08493_));
 NOR3_X1 _17774_ (.A1(_08437_),
    .A2(_08477_),
    .A3(_08493_),
    .ZN(_08494_));
 NOR3_X2 _17775_ (.A1(_08458_),
    .A2(_08491_),
    .A3(_08494_),
    .ZN(_08495_));
 OAI22_X4 _17776_ (.A1(_08439_),
    .A2(_08442_),
    .B1(_06647_),
    .B2(_06661_),
    .ZN(_08496_));
 NOR2_X2 _17777_ (.A1(_08490_),
    .A2(_08496_),
    .ZN(_08497_));
 AOI221_X2 _17778_ (.A(_06661_),
    .B1(_06641_),
    .B2(_06629_),
    .C1(_06279_),
    .C2(_06646_),
    .ZN(_08498_));
 OR2_X2 _17779_ (.A1(_08467_),
    .A2(_08498_),
    .ZN(_08499_));
 AOI221_X2 _17780_ (.A(_08497_),
    .B1(_08499_),
    .B2(net789),
    .C1(_08443_),
    .C2(net1002),
    .ZN(_08500_));
 BUF_X4 _17781_ (.A(_06692_),
    .Z(_08501_));
 AOI211_X2 _17782_ (.A(_06679_),
    .B(_08495_),
    .C1(_08500_),
    .C2(_08501_),
    .ZN(_08502_));
 INV_X8 _17783_ (.A(_08455_),
    .ZN(_08503_));
 NAND3_X1 _17784_ (.A1(_08482_),
    .A2(_08480_),
    .A3(_06692_),
    .ZN(_08504_));
 AOI221_X2 _17785_ (.A(_08448_),
    .B1(_06625_),
    .B2(_06613_),
    .C1(_06401_),
    .C2(_06646_),
    .ZN(_08505_));
 AOI21_X4 _17786_ (.A(_08455_),
    .B1(_08461_),
    .B2(_08465_),
    .ZN(_08506_));
 AOI21_X1 _17787_ (.A(_08505_),
    .B1(_08506_),
    .B2(_08458_),
    .ZN(_08507_));
 BUF_X4 _17788_ (.A(_08438_),
    .Z(_08508_));
 OAI22_X1 _17789_ (.A1(_08503_),
    .A2(_08504_),
    .B1(_08507_),
    .B2(_08508_),
    .ZN(_08509_));
 NOR2_X1 _17790_ (.A1(_08467_),
    .A2(_08498_),
    .ZN(_08510_));
 XNOR2_X2 _17791_ (.A(_08435_),
    .B(_08479_),
    .ZN(_08511_));
 MUX2_X1 _17792_ (.A(_08510_),
    .B(_08511_),
    .S(_14766_),
    .Z(_08512_));
 CLKBUF_X3 _17793_ (.A(_06695_),
    .Z(_08513_));
 AOI21_X1 _17794_ (.A(_08509_),
    .B1(_08512_),
    .B2(_08513_),
    .ZN(_08514_));
 AOI21_X1 _17795_ (.A(_08502_),
    .B1(_08514_),
    .B2(_00396_),
    .ZN(_08515_));
 CLKBUF_X3 _17796_ (.A(_06716_),
    .Z(_08516_));
 MUX2_X1 _17797_ (.A(_08488_),
    .B(_08515_),
    .S(_08516_),
    .Z(_08517_));
 CLKBUF_X3 _17798_ (.A(_08459_),
    .Z(_08518_));
 CLKBUF_X3 _17799_ (.A(_08436_),
    .Z(_08519_));
 BUF_X4 _17800_ (.A(_14769_),
    .Z(_08520_));
 CLKBUF_X3 _17801_ (.A(_08461_),
    .Z(_08521_));
 CLKBUF_X3 _17802_ (.A(_08465_),
    .Z(_08522_));
 AOI21_X1 _17803_ (.A(_08520_),
    .B1(_08521_),
    .B2(_08522_),
    .ZN(_08523_));
 NOR3_X2 _17804_ (.A1(_08446_),
    .A2(_08447_),
    .A3(_08449_),
    .ZN(_08524_));
 OAI21_X1 _17805_ (.A(_08519_),
    .B1(_08523_),
    .B2(_08524_),
    .ZN(_08525_));
 NAND2_X4 _17806_ (.A1(_08474_),
    .A2(_06662_),
    .ZN(_08526_));
 INV_X4 _17807_ (.A(net789),
    .ZN(_08527_));
 OAI21_X1 _17808_ (.A(_08525_),
    .B1(_08526_),
    .B2(_08527_),
    .ZN(_08528_));
 NAND2_X1 _17809_ (.A1(_00396_),
    .A2(_08528_),
    .ZN(_08529_));
 BUF_X4 _17810_ (.A(_08486_),
    .Z(_08530_));
 BUF_X4 _17811_ (.A(_08530_),
    .Z(_08531_));
 BUF_X4 _17812_ (.A(_06663_),
    .Z(_08532_));
 NAND2_X2 _17813_ (.A1(_06611_),
    .A2(_08532_),
    .ZN(_08533_));
 INV_X1 _17814_ (.A(_08505_),
    .ZN(_08534_));
 AOI21_X1 _17815_ (.A(_14785_),
    .B1(_08533_),
    .B2(_08534_),
    .ZN(_08535_));
 CLKBUF_X3 _17816_ (.A(_08532_),
    .Z(_08536_));
 NOR2_X1 _17817_ (.A1(_08490_),
    .A2(_08536_),
    .ZN(_08537_));
 NOR3_X1 _17818_ (.A1(_14780_),
    .A2(_08489_),
    .A3(_08537_),
    .ZN(_08538_));
 OAI21_X1 _17819_ (.A(_08531_),
    .B1(_08535_),
    .B2(_08538_),
    .ZN(_08539_));
 AOI21_X1 _17820_ (.A(_08518_),
    .B1(_08529_),
    .B2(_08539_),
    .ZN(_08540_));
 BUF_X4 _17821_ (.A(_08492_),
    .Z(_08541_));
 MUX2_X1 _17822_ (.A(_08541_),
    .B(_06611_),
    .S(_08474_),
    .Z(_08542_));
 BUF_X4 _17823_ (.A(_08479_),
    .Z(_08543_));
 OAI21_X2 _17824_ (.A(_08486_),
    .B1(_08542_),
    .B2(_08543_),
    .ZN(_08544_));
 AOI21_X1 _17825_ (.A(_06664_),
    .B1(_08519_),
    .B2(_08468_),
    .ZN(_08545_));
 OAI21_X1 _17826_ (.A(_06680_),
    .B1(_08497_),
    .B2(_08545_),
    .ZN(_08546_));
 BUF_X4 _17827_ (.A(_08443_),
    .Z(_08547_));
 AOI221_X2 _17828_ (.A(_08513_),
    .B1(_08544_),
    .B2(_08546_),
    .C1(_08547_),
    .C2(_08520_),
    .ZN(_08548_));
 CLKBUF_X3 _17829_ (.A(_08458_),
    .Z(_08549_));
 BUF_X4 _17830_ (.A(_14764_),
    .Z(_08550_));
 AOI21_X2 _17831_ (.A(_08550_),
    .B1(_08521_),
    .B2(_08522_),
    .ZN(_08551_));
 AOI221_X2 _17832_ (.A(_08551_),
    .B1(_06641_),
    .B2(_06629_),
    .C1(_06628_),
    .C2(_08480_),
    .ZN(_08552_));
 NOR2_X1 _17833_ (.A1(_06610_),
    .A2(_08479_),
    .ZN(_08553_));
 NOR2_X1 _17834_ (.A1(_08469_),
    .A2(_06664_),
    .ZN(_08554_));
 NOR3_X1 _17835_ (.A1(_08508_),
    .A2(_08553_),
    .A3(_08554_),
    .ZN(_08555_));
 OAI21_X1 _17836_ (.A(_08549_),
    .B1(_08552_),
    .B2(_08555_),
    .ZN(_08556_));
 NOR4_X4 _17837_ (.A1(_06597_),
    .A2(net542),
    .A3(_06647_),
    .A4(_06661_),
    .ZN(_08557_));
 OAI21_X1 _17838_ (.A(_08519_),
    .B1(_08557_),
    .B2(_08506_),
    .ZN(_08558_));
 CLKBUF_X3 _17839_ (.A(_08474_),
    .Z(_08559_));
 CLKBUF_X3 _17840_ (.A(_08559_),
    .Z(_08560_));
 OAI21_X1 _17841_ (.A(_08560_),
    .B1(_08551_),
    .B2(_08554_),
    .ZN(_08561_));
 NAND3_X1 _17842_ (.A1(_08513_),
    .A2(_08558_),
    .A3(_08561_),
    .ZN(_08562_));
 AND3_X1 _17843_ (.A1(_06681_),
    .A2(_08556_),
    .A3(_08562_),
    .ZN(_08563_));
 NAND2_X1 _17844_ (.A1(_06677_),
    .A2(_06693_),
    .ZN(_08564_));
 AOI21_X1 _17845_ (.A(_08469_),
    .B1(_08521_),
    .B2(_08522_),
    .ZN(_08565_));
 OAI21_X1 _17846_ (.A(_14785_),
    .B1(_08557_),
    .B2(_08565_),
    .ZN(_08566_));
 BUF_X4 _17847_ (.A(_08496_),
    .Z(_08567_));
 OR2_X1 _17848_ (.A1(_08520_),
    .A2(_08567_),
    .ZN(_08568_));
 AOI21_X1 _17849_ (.A(_08564_),
    .B1(_08566_),
    .B2(_08568_),
    .ZN(_08569_));
 CLKBUF_X3 _17850_ (.A(_08474_),
    .Z(_08570_));
 CLKBUF_X3 _17851_ (.A(_08570_),
    .Z(_08571_));
 NAND2_X1 _17852_ (.A1(_14760_),
    .A2(_08571_),
    .ZN(_08572_));
 INV_X1 _17853_ (.A(_08446_),
    .ZN(_08573_));
 AOI21_X2 _17854_ (.A(_08532_),
    .B1(_08482_),
    .B2(_08573_),
    .ZN(_08574_));
 NAND2_X1 _17855_ (.A1(_08572_),
    .A2(_08574_),
    .ZN(_08575_));
 NAND2_X1 _17856_ (.A1(_08518_),
    .A2(_08575_),
    .ZN(_08576_));
 OAI21_X1 _17857_ (.A(_06716_),
    .B1(_08544_),
    .B2(_08576_),
    .ZN(_08577_));
 OAI33_X1 _17858_ (.A1(_08516_),
    .A2(_08540_),
    .A3(_08548_),
    .B1(_08563_),
    .B2(_08569_),
    .B3(_08577_),
    .ZN(_08578_));
 MUX2_X1 _17859_ (.A(_08517_),
    .B(_08578_),
    .S(_00398_),
    .Z(_00024_));
 AOI21_X1 _17860_ (.A(_08557_),
    .B1(_06663_),
    .B2(_08492_),
    .ZN(_08579_));
 NAND3_X4 _17861_ (.A1(_08527_),
    .A2(_08461_),
    .A3(_08465_),
    .ZN(_08580_));
 NAND2_X1 _17862_ (.A1(_08470_),
    .A2(_08580_),
    .ZN(_08581_));
 MUX2_X1 _17863_ (.A(_08579_),
    .B(_08581_),
    .S(_06644_),
    .Z(_08582_));
 INV_X1 _17864_ (.A(_14769_),
    .ZN(_08583_));
 AOI21_X1 _17865_ (.A(_08583_),
    .B1(_08521_),
    .B2(_08522_),
    .ZN(_08584_));
 NOR3_X1 _17866_ (.A1(_06644_),
    .A2(_08557_),
    .A3(_08584_),
    .ZN(_08585_));
 AOI21_X1 _17867_ (.A(_08585_),
    .B1(_08511_),
    .B2(_08559_),
    .ZN(_08586_));
 MUX2_X1 _17868_ (.A(_08582_),
    .B(_08586_),
    .S(_08458_),
    .Z(_08587_));
 MUX2_X1 _17869_ (.A(_08541_),
    .B(net1001),
    .S(_06644_),
    .Z(_08588_));
 NAND2_X1 _17870_ (.A1(_00395_),
    .A2(_08501_),
    .ZN(_08589_));
 OAI22_X2 _17871_ (.A1(_00395_),
    .A2(_08588_),
    .B1(_08589_),
    .B2(_14790_),
    .ZN(_08590_));
 MUX2_X1 _17872_ (.A(_08587_),
    .B(_08590_),
    .S(_08487_),
    .Z(_08591_));
 NAND2_X1 _17873_ (.A1(_08490_),
    .A2(_08474_),
    .ZN(_08592_));
 NAND2_X1 _17874_ (.A1(_08550_),
    .A2(_08437_),
    .ZN(_08593_));
 NAND3_X1 _17875_ (.A1(_06677_),
    .A2(_08592_),
    .A3(_08593_),
    .ZN(_08594_));
 AOI21_X1 _17876_ (.A(_08479_),
    .B1(_06678_),
    .B2(_14786_),
    .ZN(_08595_));
 NAND2_X1 _17877_ (.A1(_08520_),
    .A2(_06644_),
    .ZN(_08596_));
 MUX2_X1 _17878_ (.A(_08452_),
    .B(_08435_),
    .S(_06678_),
    .Z(_08597_));
 OAI21_X1 _17879_ (.A(_08596_),
    .B1(_08597_),
    .B2(_08559_),
    .ZN(_08598_));
 AOI221_X2 _17880_ (.A(_06694_),
    .B1(_08594_),
    .B2(_08595_),
    .C1(_08598_),
    .C2(_08543_),
    .ZN(_08599_));
 NAND4_X4 _17881_ (.A1(_06613_),
    .A2(net790),
    .A3(_08461_),
    .A4(_08465_),
    .ZN(_08600_));
 AOI21_X1 _17882_ (.A(_08505_),
    .B1(_08536_),
    .B2(_08469_),
    .ZN(_08601_));
 OAI221_X2 _17883_ (.A(_08530_),
    .B1(_08600_),
    .B2(_14766_),
    .C1(_08601_),
    .C2(_08508_),
    .ZN(_08602_));
 OAI21_X2 _17884_ (.A(_08490_),
    .B1(_08447_),
    .B2(_08449_),
    .ZN(_08603_));
 NAND3_X2 _17885_ (.A1(_14769_),
    .A2(_08461_),
    .A3(_08465_),
    .ZN(_08604_));
 NAND2_X1 _17886_ (.A1(_08603_),
    .A2(_08604_),
    .ZN(_08605_));
 MUX2_X1 _17887_ (.A(_08481_),
    .B(_08605_),
    .S(_08483_),
    .Z(_08606_));
 OAI21_X1 _17888_ (.A(_08602_),
    .B1(_08606_),
    .B2(_08531_),
    .ZN(_08607_));
 AOI21_X1 _17889_ (.A(_08599_),
    .B1(_08607_),
    .B2(_00397_),
    .ZN(_08608_));
 MUX2_X1 _17890_ (.A(_08591_),
    .B(_08608_),
    .S(_00399_),
    .Z(_08609_));
 INV_X2 _17891_ (.A(_14764_),
    .ZN(_08610_));
 NAND2_X2 _17892_ (.A1(_08474_),
    .A2(_06663_),
    .ZN(_08611_));
 AOI21_X1 _17893_ (.A(_08493_),
    .B1(_08532_),
    .B2(_08435_),
    .ZN(_08612_));
 OAI22_X1 _17894_ (.A1(_08610_),
    .A2(_08611_),
    .B1(_08612_),
    .B2(_08570_),
    .ZN(_08613_));
 NAND3_X4 _17895_ (.A1(_08522_),
    .A2(_08521_),
    .A3(net789),
    .ZN(_08614_));
 NAND3_X1 _17896_ (.A1(_08482_),
    .A2(_08603_),
    .A3(_08614_),
    .ZN(_08615_));
 OR2_X1 _17897_ (.A1(_08523_),
    .A2(_08557_),
    .ZN(_08616_));
 OAI21_X1 _17898_ (.A(_08615_),
    .B1(_08616_),
    .B2(_08519_),
    .ZN(_08617_));
 MUX2_X1 _17899_ (.A(_08613_),
    .B(_08617_),
    .S(_08501_),
    .Z(_08618_));
 OAI21_X2 _17900_ (.A(_08503_),
    .B1(_06648_),
    .B2(_08448_),
    .ZN(_08619_));
 AND2_X1 _17901_ (.A1(_08619_),
    .A2(_08604_),
    .ZN(_08620_));
 OAI22_X1 _17902_ (.A1(_08541_),
    .A2(_08611_),
    .B1(_08620_),
    .B2(_08559_),
    .ZN(_08621_));
 NOR3_X1 _17903_ (.A1(net1124),
    .A2(_06626_),
    .A3(_06662_),
    .ZN(_08622_));
 AOI211_X2 _17904_ (.A(_08456_),
    .B(_08622_),
    .C1(_08499_),
    .C2(net1124),
    .ZN(_08623_));
 MUX2_X1 _17905_ (.A(_08621_),
    .B(_08623_),
    .S(_08501_),
    .Z(_08624_));
 MUX2_X1 _17906_ (.A(_08618_),
    .B(_08624_),
    .S(_08487_),
    .Z(_08625_));
 NOR3_X2 _17907_ (.A1(_08610_),
    .A2(_06648_),
    .A3(_08449_),
    .ZN(_08626_));
 NOR3_X1 _17908_ (.A1(_06644_),
    .A2(_08506_),
    .A3(_08626_),
    .ZN(_08627_));
 OAI21_X1 _17909_ (.A(_08492_),
    .B1(_08447_),
    .B2(_08449_),
    .ZN(_08628_));
 OAI21_X1 _17910_ (.A(_08628_),
    .B1(_08532_),
    .B2(_08446_),
    .ZN(_08629_));
 AOI21_X1 _17911_ (.A(_08627_),
    .B1(_08629_),
    .B2(_08559_),
    .ZN(_08630_));
 NOR3_X1 _17912_ (.A1(_08506_),
    .A2(_08557_),
    .A3(_08436_),
    .ZN(_08631_));
 OAI21_X1 _17913_ (.A(_08527_),
    .B1(_08447_),
    .B2(_08449_),
    .ZN(_08632_));
 AOI21_X1 _17914_ (.A(_08474_),
    .B1(_08632_),
    .B2(_08471_),
    .ZN(_08633_));
 OR2_X1 _17915_ (.A1(_08631_),
    .A2(_08633_),
    .ZN(_08634_));
 MUX2_X1 _17916_ (.A(_08630_),
    .B(_08634_),
    .S(_06695_),
    .Z(_08635_));
 OAI21_X1 _17917_ (.A(_08614_),
    .B1(_08480_),
    .B2(_08435_),
    .ZN(_08636_));
 AOI21_X1 _17918_ (.A(_08585_),
    .B1(_08636_),
    .B2(_06645_),
    .ZN(_08637_));
 INV_X1 _17919_ (.A(_08492_),
    .ZN(_08638_));
 OAI21_X1 _17920_ (.A(_08619_),
    .B1(_06663_),
    .B2(_08638_),
    .ZN(_08639_));
 AOI22_X1 _17921_ (.A1(_06612_),
    .A2(_08547_),
    .B1(_08639_),
    .B2(_08519_),
    .ZN(_08640_));
 MUX2_X1 _17922_ (.A(_08637_),
    .B(_08640_),
    .S(_08501_),
    .Z(_08641_));
 MUX2_X1 _17923_ (.A(_08635_),
    .B(_08641_),
    .S(_08487_),
    .Z(_08642_));
 MUX2_X1 _17924_ (.A(_08625_),
    .B(_08642_),
    .S(_08516_),
    .Z(_08643_));
 MUX2_X1 _17925_ (.A(_08609_),
    .B(_08643_),
    .S(_00398_),
    .Z(_00025_));
 OAI22_X4 _17926_ (.A1(_06597_),
    .A2(net543),
    .B1(_06648_),
    .B2(_08448_),
    .ZN(_08644_));
 NAND3_X4 _17927_ (.A1(_08490_),
    .A2(_08461_),
    .A3(_08465_),
    .ZN(_08645_));
 AOI21_X1 _17928_ (.A(_08474_),
    .B1(_08644_),
    .B2(_08645_),
    .ZN(_08646_));
 AOI21_X1 _17929_ (.A(_08482_),
    .B1(_08600_),
    .B2(_08450_),
    .ZN(_08647_));
 NOR3_X1 _17930_ (.A1(_08458_),
    .A2(_08646_),
    .A3(_08647_),
    .ZN(_08648_));
 NOR3_X2 _17931_ (.A1(_08550_),
    .A2(_06648_),
    .A3(_08448_),
    .ZN(_08649_));
 OR2_X1 _17932_ (.A1(_08565_),
    .A2(_08649_),
    .ZN(_08650_));
 AND2_X1 _17933_ (.A1(_06401_),
    .A2(net80),
    .ZN(_08651_));
 NOR2_X1 _17934_ (.A1(_06279_),
    .A2(_06617_),
    .ZN(_08652_));
 NOR2_X1 _17935_ (.A1(_06279_),
    .A2(_06615_),
    .ZN(_08653_));
 MUX2_X2 _17936_ (.A(_08652_),
    .B(_08653_),
    .S(_06624_),
    .Z(_08654_));
 OAI22_X4 _17937_ (.A1(_08651_),
    .A2(_08654_),
    .B1(_06648_),
    .B2(_08448_),
    .ZN(_08655_));
 OAI21_X1 _17938_ (.A(_08655_),
    .B1(_08532_),
    .B2(_08520_),
    .ZN(_08656_));
 MUX2_X1 _17939_ (.A(_08650_),
    .B(_08656_),
    .S(_08519_),
    .Z(_08657_));
 AOI211_X2 _17940_ (.A(_08530_),
    .B(_08648_),
    .C1(_08657_),
    .C2(_08459_),
    .ZN(_08658_));
 NOR3_X2 _17941_ (.A1(_08520_),
    .A2(_08439_),
    .A3(_08442_),
    .ZN(_08659_));
 AOI21_X4 _17942_ (.A(_08659_),
    .B1(_08452_),
    .B2(_08519_),
    .ZN(_08660_));
 OAI21_X4 _17943_ (.A(_08486_),
    .B1(_08543_),
    .B2(_08660_),
    .ZN(_08661_));
 OAI21_X1 _17944_ (.A(_08543_),
    .B1(_06645_),
    .B2(_14771_),
    .ZN(_08662_));
 AOI21_X1 _17945_ (.A(_08662_),
    .B1(_08560_),
    .B2(_08490_),
    .ZN(_08663_));
 NAND3_X4 _17946_ (.A1(_08452_),
    .A2(_08521_),
    .A3(_08522_),
    .ZN(_08664_));
 AOI21_X1 _17947_ (.A(_08483_),
    .B1(_08664_),
    .B2(_08628_),
    .ZN(_08665_));
 NOR2_X1 _17948_ (.A1(_08550_),
    .A2(_08496_),
    .ZN(_08666_));
 OAI33_X1 _17949_ (.A1(_00397_),
    .A2(_08661_),
    .A3(_08663_),
    .B1(_08665_),
    .B2(_08666_),
    .B3(_08564_),
    .ZN(_08667_));
 NOR3_X1 _17950_ (.A1(_00399_),
    .A2(_08658_),
    .A3(_08667_),
    .ZN(_08668_));
 NAND2_X1 _17951_ (.A1(_08603_),
    .A2(_08580_),
    .ZN(_08669_));
 AOI221_X2 _17952_ (.A(_08501_),
    .B1(_08467_),
    .B2(_08520_),
    .C1(_08669_),
    .C2(_08483_),
    .ZN(_08670_));
 AOI22_X1 _17953_ (.A1(_14781_),
    .A2(_00395_),
    .B1(_08547_),
    .B2(net57),
    .ZN(_08671_));
 NOR2_X1 _17954_ (.A1(_00397_),
    .A2(_08671_),
    .ZN(_08672_));
 OAI21_X1 _17955_ (.A(_08531_),
    .B1(_08670_),
    .B2(_08672_),
    .ZN(_08673_));
 NOR2_X1 _17956_ (.A1(net1124),
    .A2(_08567_),
    .ZN(_08674_));
 AOI221_X2 _17957_ (.A(_08674_),
    .B1(_08547_),
    .B2(net1002),
    .C1(_08541_),
    .C2(_08499_),
    .ZN(_08675_));
 MUX2_X1 _17958_ (.A(_08469_),
    .B(_06628_),
    .S(_08437_),
    .Z(_08676_));
 MUX2_X1 _17959_ (.A(_14788_),
    .B(_08676_),
    .S(_08536_),
    .Z(_08677_));
 MUX2_X1 _17960_ (.A(_08675_),
    .B(_08677_),
    .S(_08549_),
    .Z(_08678_));
 OAI21_X2 _17961_ (.A(_08673_),
    .B1(_08678_),
    .B2(_08531_),
    .ZN(_08679_));
 AOI21_X1 _17962_ (.A(_08668_),
    .B1(_08679_),
    .B2(_00399_),
    .ZN(_08680_));
 NAND2_X1 _17963_ (.A1(_08520_),
    .A2(_06663_),
    .ZN(_08681_));
 NAND3_X1 _17964_ (.A1(_08550_),
    .A2(_08521_),
    .A3(_08522_),
    .ZN(_08682_));
 NAND3_X1 _17965_ (.A1(_08560_),
    .A2(_08681_),
    .A3(_08682_),
    .ZN(_08683_));
 NAND3_X1 _17966_ (.A1(_08468_),
    .A2(_08521_),
    .A3(_08522_),
    .ZN(_08684_));
 AND2_X1 _17967_ (.A1(_08438_),
    .A2(_08684_),
    .ZN(_08685_));
 NAND2_X1 _17968_ (.A1(_08644_),
    .A2(_08685_),
    .ZN(_08686_));
 NAND4_X1 _17969_ (.A1(_06681_),
    .A2(_08549_),
    .A3(_08683_),
    .A4(_08686_),
    .ZN(_08687_));
 NOR2_X2 _17970_ (.A1(_06628_),
    .A2(_08479_),
    .ZN(_08688_));
 NOR3_X1 _17971_ (.A1(_08483_),
    .A2(_08688_),
    .A3(_08649_),
    .ZN(_08689_));
 INV_X2 _17972_ (.A(_14774_),
    .ZN(_08690_));
 AOI21_X1 _17973_ (.A(_08557_),
    .B1(_00395_),
    .B2(_08690_),
    .ZN(_08691_));
 AOI21_X1 _17974_ (.A(_08689_),
    .B1(_08691_),
    .B2(_14780_),
    .ZN(_08692_));
 NAND2_X1 _17975_ (.A1(_06679_),
    .A2(_06694_),
    .ZN(_08693_));
 NAND3_X1 _17976_ (.A1(_06645_),
    .A2(_08619_),
    .A3(_08684_),
    .ZN(_08694_));
 AND3_X1 _17977_ (.A1(_06695_),
    .A2(_08558_),
    .A3(_08694_),
    .ZN(_08695_));
 AOI21_X1 _17978_ (.A(_08659_),
    .B1(_08685_),
    .B2(_08655_),
    .ZN(_08696_));
 AOI21_X1 _17979_ (.A(_08695_),
    .B1(_08696_),
    .B2(_08549_),
    .ZN(_08697_));
 OAI221_X1 _17980_ (.A(_08687_),
    .B1(_08692_),
    .B2(_08693_),
    .C1(_08697_),
    .C2(_00396_),
    .ZN(_08698_));
 NAND3_X1 _17981_ (.A1(_06645_),
    .A2(_08603_),
    .A3(_08580_),
    .ZN(_08699_));
 OR3_X1 _17982_ (.A1(_08570_),
    .A2(_08505_),
    .A3(_08489_),
    .ZN(_08700_));
 NAND3_X1 _17983_ (.A1(_08501_),
    .A2(_08699_),
    .A3(_08700_),
    .ZN(_08701_));
 MUX2_X1 _17984_ (.A(_08467_),
    .B(_08498_),
    .S(_06627_),
    .Z(_08702_));
 OAI21_X1 _17985_ (.A(_08655_),
    .B1(_08474_),
    .B2(_06626_),
    .ZN(_08703_));
 OAI21_X1 _17986_ (.A(_08600_),
    .B1(_08436_),
    .B2(_06628_),
    .ZN(_08704_));
 AOI221_X1 _17987_ (.A(_08702_),
    .B1(_08703_),
    .B2(_06610_),
    .C1(_08704_),
    .C2(_08503_),
    .ZN(_08705_));
 OAI21_X1 _17988_ (.A(_08701_),
    .B1(_08705_),
    .B2(_08459_),
    .ZN(_08706_));
 NAND2_X1 _17989_ (.A1(_08503_),
    .A2(_06643_),
    .ZN(_08707_));
 AOI21_X1 _17990_ (.A(_06662_),
    .B1(_08436_),
    .B2(net1230),
    .ZN(_08708_));
 AOI221_X2 _17991_ (.A(_06692_),
    .B1(_08708_),
    .B2(_08707_),
    .C1(_08480_),
    .C2(_14783_),
    .ZN(_08709_));
 MUX2_X1 _17992_ (.A(_06611_),
    .B(_08436_),
    .S(_08435_),
    .Z(_08710_));
 MUX2_X1 _17993_ (.A(_14790_),
    .B(_08710_),
    .S(_06664_),
    .Z(_08711_));
 AOI21_X1 _17994_ (.A(_08709_),
    .B1(_08711_),
    .B2(_08549_),
    .ZN(_08712_));
 MUX2_X1 _17995_ (.A(_08706_),
    .B(_08712_),
    .S(_08487_),
    .Z(_08713_));
 MUX2_X1 _17996_ (.A(_08698_),
    .B(_08713_),
    .S(_00399_),
    .Z(_08714_));
 MUX2_X1 _17997_ (.A(_08680_),
    .B(_08714_),
    .S(_00398_),
    .Z(_00026_));
 AOI21_X1 _17998_ (.A(_08557_),
    .B1(_08482_),
    .B2(net992),
    .ZN(_08715_));
 AOI221_X2 _17999_ (.A(_06694_),
    .B1(_08547_),
    .B2(_14761_),
    .C1(_08715_),
    .C2(_08550_),
    .ZN(_08716_));
 AOI221_X2 _18000_ (.A(_08458_),
    .B1(_08498_),
    .B2(net992),
    .C1(_08510_),
    .C2(_08468_),
    .ZN(_08717_));
 NAND3_X1 _18001_ (.A1(_08503_),
    .A2(_08521_),
    .A3(_08522_),
    .ZN(_08718_));
 NAND2_X1 _18002_ (.A1(net1235),
    .A2(_06695_),
    .ZN(_08719_));
 NAND3_X1 _18003_ (.A1(_08644_),
    .A2(_08718_),
    .A3(_08719_),
    .ZN(_08720_));
 OAI221_X1 _18004_ (.A(_08531_),
    .B1(_08716_),
    .B2(_08717_),
    .C1(_08720_),
    .C2(_14785_),
    .ZN(_08721_));
 NAND2_X1 _18005_ (.A1(_14771_),
    .A2(_08498_),
    .ZN(_08722_));
 NOR3_X4 _18006_ (.A1(net1001),
    .A2(_06648_),
    .A3(_08448_),
    .ZN(_08723_));
 OAI21_X1 _18007_ (.A(_06645_),
    .B1(_08506_),
    .B2(_08723_),
    .ZN(_08724_));
 AOI21_X1 _18008_ (.A(_06695_),
    .B1(_08722_),
    .B2(_08724_),
    .ZN(_08725_));
 NAND3_X1 _18009_ (.A1(_08503_),
    .A2(_08543_),
    .A3(_06694_),
    .ZN(_08726_));
 AOI21_X1 _18010_ (.A(_08560_),
    .B1(_08450_),
    .B2(_08726_),
    .ZN(_08727_));
 OR3_X1 _18011_ (.A1(_08487_),
    .A2(_08725_),
    .A3(_08727_),
    .ZN(_08728_));
 AOI21_X1 _18012_ (.A(_00399_),
    .B1(_08721_),
    .B2(_08728_),
    .ZN(_08729_));
 NAND2_X1 _18013_ (.A1(_08482_),
    .A2(_06678_),
    .ZN(_08730_));
 NAND3_X1 _18014_ (.A1(_08570_),
    .A2(_08480_),
    .A3(_06677_),
    .ZN(_08731_));
 AOI21_X1 _18015_ (.A(net1235),
    .B1(_08730_),
    .B2(_08731_),
    .ZN(_08732_));
 OAI21_X1 _18016_ (.A(_08490_),
    .B1(_08483_),
    .B2(_06680_),
    .ZN(_08733_));
 NAND3_X1 _18017_ (.A1(_14760_),
    .A2(_08571_),
    .A3(_08486_),
    .ZN(_08734_));
 NAND4_X1 _18018_ (.A1(_00395_),
    .A2(_08730_),
    .A3(_08733_),
    .A4(_08734_),
    .ZN(_08735_));
 CLKBUF_X3 _18019_ (.A(_08543_),
    .Z(_08736_));
 NAND3_X1 _18020_ (.A1(_14760_),
    .A2(_08571_),
    .A3(_06680_),
    .ZN(_08737_));
 NAND3_X1 _18021_ (.A1(net1235),
    .A2(_14771_),
    .A3(_08530_),
    .ZN(_08738_));
 NAND3_X1 _18022_ (.A1(_08736_),
    .A2(_08737_),
    .A3(_08738_),
    .ZN(_08739_));
 AOI21_X1 _18023_ (.A(_08732_),
    .B1(_08735_),
    .B2(_08739_),
    .ZN(_08740_));
 OAI221_X1 _18024_ (.A(_08645_),
    .B1(_08442_),
    .B2(_08439_),
    .C1(_08550_),
    .C2(_08543_),
    .ZN(_08741_));
 OAI21_X1 _18025_ (.A(_08583_),
    .B1(_08447_),
    .B2(_08449_),
    .ZN(_08742_));
 NAND3_X1 _18026_ (.A1(_08560_),
    .A2(_08600_),
    .A3(_08742_),
    .ZN(_08743_));
 NAND3_X1 _18027_ (.A1(_08487_),
    .A2(_08741_),
    .A3(_08743_),
    .ZN(_08744_));
 NOR3_X1 _18028_ (.A1(_08571_),
    .A2(_08477_),
    .A3(_08723_),
    .ZN(_08745_));
 AOI21_X1 _18029_ (.A(_08506_),
    .B1(_08736_),
    .B2(_14761_),
    .ZN(_08746_));
 AOI21_X1 _18030_ (.A(_08745_),
    .B1(_08746_),
    .B2(_14785_),
    .ZN(_08747_));
 OAI21_X1 _18031_ (.A(_08744_),
    .B1(_08747_),
    .B2(_08531_),
    .ZN(_08748_));
 MUX2_X1 _18032_ (.A(_08740_),
    .B(_08748_),
    .S(_00397_),
    .Z(_08749_));
 AOI21_X1 _18033_ (.A(_08729_),
    .B1(_08749_),
    .B2(_00399_),
    .ZN(_08750_));
 NAND2_X1 _18034_ (.A1(_06664_),
    .A2(_06694_),
    .ZN(_08751_));
 OAI221_X1 _18035_ (.A(_08571_),
    .B1(_08536_),
    .B2(_08550_),
    .C1(_08751_),
    .C2(net1235),
    .ZN(_08752_));
 NAND3_X1 _18036_ (.A1(net1116),
    .A2(_08543_),
    .A3(_08458_),
    .ZN(_08753_));
 OAI21_X2 _18037_ (.A(_08468_),
    .B1(_08447_),
    .B2(_08449_),
    .ZN(_08754_));
 NAND2_X2 _18038_ (.A1(_08645_),
    .A2(_08754_),
    .ZN(_08755_));
 OAI21_X1 _18039_ (.A(_08753_),
    .B1(_08755_),
    .B2(_08501_),
    .ZN(_08756_));
 OAI21_X1 _18040_ (.A(_08752_),
    .B1(_08756_),
    .B2(_14785_),
    .ZN(_08757_));
 AND2_X1 _18041_ (.A1(_08436_),
    .A2(_08600_),
    .ZN(_08758_));
 OAI222_X2 _18042_ (.A1(net524),
    .A2(_08567_),
    .B1(_08758_),
    .B2(_06612_),
    .C1(_06628_),
    .C2(_08526_),
    .ZN(_08759_));
 AOI21_X1 _18043_ (.A(_08690_),
    .B1(_08521_),
    .B2(_08522_),
    .ZN(_08760_));
 NOR3_X2 _18044_ (.A1(_08760_),
    .A2(_08723_),
    .A3(_08437_),
    .ZN(_08761_));
 OAI21_X2 _18045_ (.A(_08644_),
    .B1(_08532_),
    .B2(_08638_),
    .ZN(_08762_));
 AOI21_X1 _18046_ (.A(_08761_),
    .B1(_08762_),
    .B2(_08438_),
    .ZN(_08763_));
 MUX2_X1 _18047_ (.A(_08759_),
    .B(_08763_),
    .S(_08501_),
    .Z(_08764_));
 MUX2_X1 _18048_ (.A(_08757_),
    .B(_08764_),
    .S(_08487_),
    .Z(_08765_));
 MUX2_X1 _18049_ (.A(_08435_),
    .B(_08436_),
    .S(_06610_),
    .Z(_08766_));
 AOI221_X2 _18050_ (.A(_06694_),
    .B1(_08467_),
    .B2(net57),
    .C1(_08766_),
    .C2(_08480_),
    .ZN(_08767_));
 AND3_X1 _18051_ (.A1(_08570_),
    .A2(_08645_),
    .A3(_08470_),
    .ZN(_08768_));
 NOR3_X1 _18052_ (.A1(_06645_),
    .A2(_08489_),
    .A3(_08493_),
    .ZN(_08769_));
 NOR3_X1 _18053_ (.A1(_08459_),
    .A2(_08768_),
    .A3(_08769_),
    .ZN(_08770_));
 NOR3_X2 _18054_ (.A1(_08767_),
    .A2(_08770_),
    .A3(_06681_),
    .ZN(_08771_));
 AOI21_X1 _18055_ (.A(_08570_),
    .B1(_08718_),
    .B2(_08655_),
    .ZN(_08772_));
 OAI21_X1 _18056_ (.A(_08550_),
    .B1(_08447_),
    .B2(_08449_),
    .ZN(_08773_));
 AOI21_X1 _18057_ (.A(_08519_),
    .B1(_08684_),
    .B2(_08773_),
    .ZN(_08774_));
 OR3_X1 _18058_ (.A1(_06695_),
    .A2(_08772_),
    .A3(_08774_),
    .ZN(_08775_));
 AOI221_X1 _18059_ (.A(_08646_),
    .B1(_08553_),
    .B2(_06628_),
    .C1(net1002),
    .C2(_08547_),
    .ZN(_08776_));
 OAI21_X1 _18060_ (.A(_08775_),
    .B1(_08776_),
    .B2(_08518_),
    .ZN(_08777_));
 AOI21_X1 _18061_ (.A(_08771_),
    .B1(_08777_),
    .B2(_00396_),
    .ZN(_08778_));
 MUX2_X1 _18062_ (.A(_08765_),
    .B(_08778_),
    .S(_00399_),
    .Z(_08779_));
 MUX2_X1 _18063_ (.A(_08750_),
    .B(_08779_),
    .S(_00398_),
    .Z(_00027_));
 NAND2_X1 _18064_ (.A1(net992),
    .A2(_08482_),
    .ZN(_08780_));
 AOI21_X1 _18065_ (.A(_08479_),
    .B1(_08570_),
    .B2(_08690_),
    .ZN(_08781_));
 AOI21_X1 _18066_ (.A(_08486_),
    .B1(_08780_),
    .B2(_08781_),
    .ZN(_08782_));
 NAND2_X1 _18067_ (.A1(net789),
    .A2(_08570_),
    .ZN(_08783_));
 AOI21_X2 _18068_ (.A(_06679_),
    .B1(_08574_),
    .B2(_08783_),
    .ZN(_08784_));
 NAND3_X1 _18069_ (.A1(net1116),
    .A2(_14771_),
    .A3(_08536_),
    .ZN(_08785_));
 AOI21_X1 _18070_ (.A(_08782_),
    .B1(_08784_),
    .B2(_08785_),
    .ZN(_08786_));
 OAI21_X1 _18071_ (.A(_08459_),
    .B1(_08722_),
    .B2(_08784_),
    .ZN(_08787_));
 OAI22_X2 _18072_ (.A1(_06681_),
    .A2(_08567_),
    .B1(_08784_),
    .B2(_08534_),
    .ZN(_08788_));
 AOI211_X2 _18073_ (.A(_08786_),
    .B(_08787_),
    .C1(_14761_),
    .C2(_08788_),
    .ZN(_08789_));
 OAI21_X1 _18074_ (.A(_14780_),
    .B1(_08475_),
    .B2(_08688_),
    .ZN(_08790_));
 AOI21_X1 _18075_ (.A(_08487_),
    .B1(_08467_),
    .B2(_08468_),
    .ZN(_08791_));
 NAND2_X1 _18076_ (.A1(_08541_),
    .A2(_08736_),
    .ZN(_08792_));
 OAI21_X1 _18077_ (.A(_08792_),
    .B1(_08592_),
    .B2(_08736_),
    .ZN(_08793_));
 AOI22_X1 _18078_ (.A1(_08790_),
    .A2(_08791_),
    .B1(_08793_),
    .B2(_08531_),
    .ZN(_08794_));
 OAI21_X1 _18079_ (.A(_08516_),
    .B1(_08794_),
    .B2(_08518_),
    .ZN(_08795_));
 AOI21_X1 _18080_ (.A(_08459_),
    .B1(_08508_),
    .B2(_08690_),
    .ZN(_08796_));
 OAI21_X1 _18081_ (.A(_08796_),
    .B1(_08605_),
    .B2(_14780_),
    .ZN(_08797_));
 NAND3_X1 _18082_ (.A1(_08508_),
    .A2(_08470_),
    .A3(_08604_),
    .ZN(_08798_));
 NAND2_X1 _18083_ (.A1(_08655_),
    .A2(_08682_),
    .ZN(_08799_));
 OAI21_X1 _18084_ (.A(_08798_),
    .B1(_08799_),
    .B2(_14780_),
    .ZN(_08800_));
 OAI221_X1 _18085_ (.A(_08797_),
    .B1(_08800_),
    .B2(_08513_),
    .C1(_06665_),
    .C2(_06676_),
    .ZN(_08801_));
 NAND3_X1 _18086_ (.A1(_08560_),
    .A2(_08655_),
    .A3(_08604_),
    .ZN(_08802_));
 AOI21_X1 _18087_ (.A(_08513_),
    .B1(_08478_),
    .B2(_08802_),
    .ZN(_08803_));
 OAI21_X1 _18088_ (.A(_14780_),
    .B1(_08565_),
    .B2(_08649_),
    .ZN(_08804_));
 OAI21_X1 _18089_ (.A(_08804_),
    .B1(_08755_),
    .B2(_14780_),
    .ZN(_08805_));
 AOI21_X1 _18090_ (.A(_08803_),
    .B1(_08805_),
    .B2(_00397_),
    .ZN(_08806_));
 OAI21_X1 _18091_ (.A(_08801_),
    .B1(_08806_),
    .B2(_00396_),
    .ZN(_08807_));
 OAI22_X1 _18092_ (.A1(_08789_),
    .A2(_08795_),
    .B1(_08807_),
    .B2(_08516_),
    .ZN(_08808_));
 NAND3_X1 _18093_ (.A1(_08571_),
    .A2(_08655_),
    .A3(_08614_),
    .ZN(_08809_));
 NAND3_X1 _18094_ (.A1(_08530_),
    .A2(_08780_),
    .A3(_08809_),
    .ZN(_08810_));
 OAI21_X1 _18095_ (.A(_08754_),
    .B1(_08524_),
    .B2(_08560_),
    .ZN(_08811_));
 OAI21_X1 _18096_ (.A(_08810_),
    .B1(_08811_),
    .B2(_08487_),
    .ZN(_08812_));
 OAI21_X1 _18097_ (.A(_08707_),
    .B1(_14785_),
    .B2(_08583_),
    .ZN(_08813_));
 AOI21_X1 _18098_ (.A(_08544_),
    .B1(_08813_),
    .B2(_08736_),
    .ZN(_08814_));
 NAND3_X1 _18099_ (.A1(_14785_),
    .A2(_06680_),
    .A3(_08629_),
    .ZN(_08815_));
 NAND2_X1 _18100_ (.A1(_06716_),
    .A2(_08815_),
    .ZN(_08816_));
 OAI22_X1 _18101_ (.A1(_06716_),
    .A2(_08812_),
    .B1(_08814_),
    .B2(_08816_),
    .ZN(_08817_));
 NOR2_X1 _18102_ (.A1(_06612_),
    .A2(_08532_),
    .ZN(_08818_));
 NAND2_X1 _18103_ (.A1(_14771_),
    .A2(_08571_),
    .ZN(_08819_));
 OAI221_X2 _18104_ (.A(_06679_),
    .B1(_08611_),
    .B2(_08527_),
    .C1(_08435_),
    .C2(_06645_),
    .ZN(_08820_));
 NOR2_X1 _18105_ (.A1(_06628_),
    .A2(_08437_),
    .ZN(_08821_));
 AOI21_X1 _18106_ (.A(_08547_),
    .B1(_08482_),
    .B2(net992),
    .ZN(_08822_));
 OAI221_X2 _18107_ (.A(_08486_),
    .B1(_08533_),
    .B2(_08821_),
    .C1(_08822_),
    .C2(_14771_),
    .ZN(_08823_));
 AOI22_X2 _18108_ (.A1(_08818_),
    .A2(_08819_),
    .B1(_08820_),
    .B2(_08823_),
    .ZN(_08824_));
 NAND2_X1 _18109_ (.A1(_08437_),
    .A2(_08479_),
    .ZN(_08825_));
 OAI22_X1 _18110_ (.A1(_14761_),
    .A2(_08825_),
    .B1(_08649_),
    .B2(_08519_),
    .ZN(_08826_));
 AOI21_X2 _18111_ (.A(_06644_),
    .B1(_08614_),
    .B2(_08742_),
    .ZN(_08827_));
 AOI21_X1 _18112_ (.A(_08827_),
    .B1(_08511_),
    .B2(_06645_),
    .ZN(_08828_));
 MUX2_X1 _18113_ (.A(_08826_),
    .B(_08828_),
    .S(_06680_),
    .Z(_08829_));
 MUX2_X1 _18114_ (.A(_08824_),
    .B(_08829_),
    .S(_06716_),
    .Z(_08830_));
 MUX2_X1 _18115_ (.A(_08817_),
    .B(_08830_),
    .S(_08518_),
    .Z(_08831_));
 MUX2_X1 _18116_ (.A(_08808_),
    .B(_08831_),
    .S(_00398_),
    .Z(_00028_));
 NOR2_X1 _18117_ (.A1(_08477_),
    .A2(_08626_),
    .ZN(_08832_));
 OAI221_X1 _18118_ (.A(_08530_),
    .B1(_08567_),
    .B2(_08490_),
    .C1(_08832_),
    .C2(_08508_),
    .ZN(_08833_));
 AND2_X1 _18119_ (.A1(_08603_),
    .A2(_08471_),
    .ZN(_08834_));
 OAI221_X1 _18120_ (.A(_06680_),
    .B1(_08825_),
    .B2(_14760_),
    .C1(_08834_),
    .C2(_08508_),
    .ZN(_08835_));
 AOI21_X1 _18121_ (.A(_06716_),
    .B1(_08833_),
    .B2(_08835_),
    .ZN(_08836_));
 OAI21_X1 _18122_ (.A(_06645_),
    .B1(_08489_),
    .B2(_08626_),
    .ZN(_08837_));
 NAND3_X1 _18123_ (.A1(_08483_),
    .A2(_08645_),
    .A3(_08619_),
    .ZN(_08838_));
 AOI21_X1 _18124_ (.A(_08530_),
    .B1(_08837_),
    .B2(_08838_),
    .ZN(_08839_));
 AOI221_X2 _18125_ (.A(_06678_),
    .B1(_08498_),
    .B2(_08541_),
    .C1(net1001),
    .C2(_06664_),
    .ZN(_08840_));
 NOR3_X1 _18126_ (.A1(_06717_),
    .A2(_08839_),
    .A3(_08840_),
    .ZN(_08841_));
 OR3_X1 _18127_ (.A1(_00397_),
    .A2(_08836_),
    .A3(_08841_),
    .ZN(_08842_));
 NAND2_X1 _18128_ (.A1(_08536_),
    .A2(_06679_),
    .ZN(_08843_));
 AOI21_X1 _18129_ (.A(_08547_),
    .B1(_08486_),
    .B2(_08435_),
    .ZN(_08844_));
 OAI222_X2 _18130_ (.A1(_14760_),
    .A2(_08731_),
    .B1(_08843_),
    .B2(_08588_),
    .C1(_08844_),
    .C2(_14761_),
    .ZN(_08845_));
 MUX2_X1 _18131_ (.A(_08536_),
    .B(_08818_),
    .S(_06680_),
    .Z(_08846_));
 AOI21_X1 _18132_ (.A(_08845_),
    .B1(_08846_),
    .B2(_14760_),
    .ZN(_08847_));
 AOI221_X2 _18133_ (.A(_06679_),
    .B1(_08547_),
    .B2(net57),
    .C1(_08762_),
    .C2(_08519_),
    .ZN(_08848_));
 AOI22_X1 _18134_ (.A1(_08736_),
    .A2(_08596_),
    .B1(_08467_),
    .B2(_08610_),
    .ZN(_08849_));
 AOI21_X1 _18135_ (.A(_08848_),
    .B1(_08849_),
    .B2(_06681_),
    .ZN(_08850_));
 MUX2_X1 _18136_ (.A(_08847_),
    .B(_08850_),
    .S(_06716_),
    .Z(_08851_));
 OAI21_X1 _18137_ (.A(_08842_),
    .B1(_08851_),
    .B2(_08518_),
    .ZN(_08852_));
 AND3_X1 _18138_ (.A1(_08559_),
    .A2(_08681_),
    .A3(_08684_),
    .ZN(_08853_));
 AOI21_X4 _18139_ (.A(_08559_),
    .B1(_08644_),
    .B2(_08664_),
    .ZN(_08854_));
 OAI21_X2 _18140_ (.A(_06695_),
    .B1(_08854_),
    .B2(_08853_),
    .ZN(_08855_));
 OAI21_X4 _18141_ (.A(net1230),
    .B1(_08447_),
    .B2(_08448_),
    .ZN(_08856_));
 AOI221_X2 _18142_ (.A(_06693_),
    .B1(_06643_),
    .B2(_08856_),
    .C1(_08479_),
    .C2(_08520_),
    .ZN(_08857_));
 NOR2_X2 _18143_ (.A1(_08857_),
    .A2(_08530_),
    .ZN(_08858_));
 OAI21_X1 _18144_ (.A(_08559_),
    .B1(_08505_),
    .B2(_08551_),
    .ZN(_08859_));
 AOI21_X1 _18145_ (.A(_08458_),
    .B1(_08525_),
    .B2(_08859_),
    .ZN(_08860_));
 NAND3_X1 _18146_ (.A1(_08438_),
    .A2(_08645_),
    .A3(_08754_),
    .ZN(_08861_));
 OAI21_X1 _18147_ (.A(_08861_),
    .B1(_08644_),
    .B2(_08483_),
    .ZN(_08862_));
 AOI21_X1 _18148_ (.A(_08860_),
    .B1(_08862_),
    .B2(_08459_),
    .ZN(_08863_));
 AOI221_X2 _18149_ (.A(_06716_),
    .B1(_08855_),
    .B2(_08858_),
    .C1(_08863_),
    .C2(_08531_),
    .ZN(_08864_));
 NOR4_X1 _18150_ (.A1(_14761_),
    .A2(_06628_),
    .A3(_08532_),
    .A4(_06692_),
    .ZN(_08865_));
 OAI22_X1 _18151_ (.A1(_08583_),
    .A2(_08526_),
    .B1(_08567_),
    .B2(_08541_),
    .ZN(_08866_));
 OAI21_X1 _18152_ (.A(_08570_),
    .B1(_08532_),
    .B2(_06694_),
    .ZN(_08867_));
 NAND3_X1 _18153_ (.A1(_08504_),
    .A2(_08751_),
    .A3(_08867_),
    .ZN(_08868_));
 AOI221_X1 _18154_ (.A(_08865_),
    .B1(_08866_),
    .B2(_08458_),
    .C1(_08868_),
    .C2(_14761_),
    .ZN(_08869_));
 NAND2_X1 _18155_ (.A1(_08638_),
    .A2(_08498_),
    .ZN(_08870_));
 NAND3_X1 _18156_ (.A1(_08549_),
    .A2(_08870_),
    .A3(_08837_),
    .ZN(_08871_));
 NAND3_X1 _18157_ (.A1(_08508_),
    .A2(_08600_),
    .A3(_08619_),
    .ZN(_08872_));
 OAI21_X1 _18158_ (.A(_08856_),
    .B1(_00395_),
    .B2(_08468_),
    .ZN(_08873_));
 OAI21_X1 _18159_ (.A(_08872_),
    .B1(_08873_),
    .B2(_14780_),
    .ZN(_08874_));
 OAI21_X1 _18160_ (.A(_08871_),
    .B1(_08874_),
    .B2(_08518_),
    .ZN(_08875_));
 MUX2_X1 _18161_ (.A(_08869_),
    .B(_08875_),
    .S(_00396_),
    .Z(_08876_));
 AOI21_X1 _18162_ (.A(_08864_),
    .B1(_08876_),
    .B2(_08516_),
    .ZN(_08877_));
 MUX2_X1 _18163_ (.A(_08852_),
    .B(_08877_),
    .S(_00398_),
    .Z(_00029_));
 INV_X1 _18164_ (.A(_14782_),
    .ZN(_08878_));
 MUX2_X1 _18165_ (.A(_08690_),
    .B(_06627_),
    .S(_08436_),
    .Z(_08879_));
 MUX2_X1 _18166_ (.A(_08878_),
    .B(_08879_),
    .S(_08480_),
    .Z(_08880_));
 NOR2_X1 _18167_ (.A1(_08486_),
    .A2(_08497_),
    .ZN(_08881_));
 NOR2_X1 _18168_ (.A1(_08610_),
    .A2(_08480_),
    .ZN(_08882_));
 OAI21_X1 _18169_ (.A(_08571_),
    .B1(_08818_),
    .B2(_08882_),
    .ZN(_08883_));
 AOI22_X1 _18170_ (.A1(_08530_),
    .A2(_08880_),
    .B1(_08881_),
    .B2(_08883_),
    .ZN(_08884_));
 OAI21_X1 _18171_ (.A(_06680_),
    .B1(_08567_),
    .B2(_14760_),
    .ZN(_08885_));
 OAI21_X2 _18172_ (.A(_08661_),
    .B1(_08761_),
    .B2(_08885_),
    .ZN(_08886_));
 MUX2_X1 _18173_ (.A(_08884_),
    .B(_08886_),
    .S(_08549_),
    .Z(_08887_));
 NOR2_X1 _18174_ (.A1(net57),
    .A2(_08567_),
    .ZN(_08888_));
 AOI21_X1 _18175_ (.A(_08723_),
    .B1(_08536_),
    .B2(_14771_),
    .ZN(_08889_));
 NOR3_X1 _18176_ (.A1(_08508_),
    .A2(_08530_),
    .A3(_08889_),
    .ZN(_08890_));
 OAI21_X1 _18177_ (.A(_08549_),
    .B1(_08888_),
    .B2(_08890_),
    .ZN(_08891_));
 MUX2_X1 _18178_ (.A(_08503_),
    .B(_08452_),
    .S(_06644_),
    .Z(_08892_));
 MUX2_X1 _18179_ (.A(_14781_),
    .B(_08892_),
    .S(_08736_),
    .Z(_08893_));
 AOI22_X1 _18180_ (.A1(_08503_),
    .A2(_08547_),
    .B1(_08499_),
    .B2(_06612_),
    .ZN(_08894_));
 AOI21_X1 _18181_ (.A(_08772_),
    .B1(_08472_),
    .B2(_08571_),
    .ZN(_08895_));
 MUX2_X1 _18182_ (.A(_08894_),
    .B(_08895_),
    .S(_06695_),
    .Z(_08896_));
 OAI221_X1 _18183_ (.A(_08891_),
    .B1(_08893_),
    .B2(_08693_),
    .C1(_08896_),
    .C2(_06681_),
    .ZN(_08897_));
 MUX2_X1 _18184_ (.A(_08887_),
    .B(_08897_),
    .S(_00399_),
    .Z(_08898_));
 MUX2_X1 _18185_ (.A(net57),
    .B(net1116),
    .S(_08482_),
    .Z(_08899_));
 MUX2_X1 _18186_ (.A(_14786_),
    .B(_08899_),
    .S(_08736_),
    .Z(_08900_));
 OAI22_X1 _18187_ (.A1(net1235),
    .A2(_14780_),
    .B1(_08825_),
    .B2(_08550_),
    .ZN(_08901_));
 NAND2_X1 _18188_ (.A1(_00397_),
    .A2(_08785_),
    .ZN(_08902_));
 OAI221_X1 _18189_ (.A(_00396_),
    .B1(_00397_),
    .B2(_08900_),
    .C1(_08901_),
    .C2(_08902_),
    .ZN(_08903_));
 AOI21_X1 _18190_ (.A(_08438_),
    .B1(_06664_),
    .B2(net1116),
    .ZN(_08904_));
 OAI222_X2 _18191_ (.A1(_08469_),
    .A2(_08526_),
    .B1(_08567_),
    .B2(net1235),
    .C1(_08904_),
    .C2(_14771_),
    .ZN(_08905_));
 OR2_X1 _18192_ (.A1(_08513_),
    .A2(_08904_),
    .ZN(_08906_));
 NOR2_X1 _18193_ (.A1(_14785_),
    .A2(_08755_),
    .ZN(_08907_));
 OAI221_X1 _18194_ (.A(_08531_),
    .B1(_08518_),
    .B2(_08905_),
    .C1(_08906_),
    .C2(_08907_),
    .ZN(_08908_));
 NAND3_X1 _18195_ (.A1(_08516_),
    .A2(_08903_),
    .A3(_08908_),
    .ZN(_08909_));
 NAND2_X1 _18196_ (.A1(_08580_),
    .A2(_08754_),
    .ZN(_08910_));
 AOI221_X1 _18197_ (.A(_08693_),
    .B1(_08910_),
    .B2(_08438_),
    .C1(_08467_),
    .C2(_08446_),
    .ZN(_08911_));
 NOR2_X1 _18198_ (.A1(_06679_),
    .A2(_06694_),
    .ZN(_08912_));
 MUX2_X1 _18199_ (.A(_08610_),
    .B(_08690_),
    .S(_06644_),
    .Z(_08913_));
 OAI21_X1 _18200_ (.A(_08912_),
    .B1(_08913_),
    .B2(_08536_),
    .ZN(_08914_));
 NOR2_X1 _18201_ (.A1(_08638_),
    .A2(_08438_),
    .ZN(_08915_));
 AOI21_X1 _18202_ (.A(_08915_),
    .B1(_08508_),
    .B2(_08573_),
    .ZN(_08916_));
 AOI21_X1 _18203_ (.A(_08914_),
    .B1(_08916_),
    .B2(_00395_),
    .ZN(_08917_));
 AOI221_X1 _18204_ (.A(_08564_),
    .B1(_08611_),
    .B2(_06628_),
    .C1(_08688_),
    .C2(_14761_),
    .ZN(_08918_));
 NAND3_X1 _18205_ (.A1(_08468_),
    .A2(_08438_),
    .A3(_06664_),
    .ZN(_08919_));
 AND4_X1 _18206_ (.A1(_06680_),
    .A2(_08501_),
    .A3(_08894_),
    .A4(_08919_),
    .ZN(_08920_));
 OR4_X1 _18207_ (.A1(_08911_),
    .A2(_08917_),
    .A3(_08918_),
    .A4(_08920_),
    .ZN(_08921_));
 OAI21_X1 _18208_ (.A(_08909_),
    .B1(_08921_),
    .B2(_08516_),
    .ZN(_08922_));
 MUX2_X1 _18209_ (.A(_08898_),
    .B(_08922_),
    .S(_00398_),
    .Z(_00030_));
 NAND3_X1 _18210_ (.A1(net792),
    .A2(_06663_),
    .A3(_06678_),
    .ZN(_08923_));
 AOI21_X1 _18211_ (.A(_06644_),
    .B1(_08645_),
    .B2(_08923_),
    .ZN(_08924_));
 OAI21_X1 _18212_ (.A(_08526_),
    .B1(_06678_),
    .B2(_08479_),
    .ZN(_08925_));
 AOI221_X1 _18213_ (.A(_08924_),
    .B1(_06677_),
    .B2(_08570_),
    .C1(_08541_),
    .C2(_08925_),
    .ZN(_08926_));
 OR2_X1 _18214_ (.A1(_08541_),
    .A2(_08731_),
    .ZN(_08927_));
 OR2_X1 _18215_ (.A1(_08533_),
    .A2(_08730_),
    .ZN(_08928_));
 NOR3_X1 _18216_ (.A1(_08559_),
    .A2(_06664_),
    .A3(_06679_),
    .ZN(_08929_));
 OAI21_X1 _18217_ (.A(_14760_),
    .B1(_08467_),
    .B2(_08929_),
    .ZN(_08930_));
 NOR3_X1 _18218_ (.A1(_08435_),
    .A2(_08480_),
    .A3(_06679_),
    .ZN(_08931_));
 NOR2_X1 _18219_ (.A1(_06664_),
    .A2(_08486_),
    .ZN(_08932_));
 OAI21_X1 _18220_ (.A(_14761_),
    .B1(_08931_),
    .B2(_08932_),
    .ZN(_08933_));
 NAND4_X1 _18221_ (.A1(_08927_),
    .A2(_08928_),
    .A3(_08930_),
    .A4(_08933_),
    .ZN(_08934_));
 MUX2_X1 _18222_ (.A(_08926_),
    .B(_08934_),
    .S(_08513_),
    .Z(_08935_));
 AOI21_X2 _18223_ (.A(_08559_),
    .B1(_08664_),
    .B2(_08742_),
    .ZN(_08936_));
 AOI21_X1 _18224_ (.A(_08936_),
    .B1(_08511_),
    .B2(_08571_),
    .ZN(_08937_));
 AOI21_X1 _18225_ (.A(_06694_),
    .B1(_08543_),
    .B2(_14783_),
    .ZN(_08938_));
 OAI21_X1 _18226_ (.A(_08938_),
    .B1(_08567_),
    .B2(_08490_),
    .ZN(_08939_));
 OAI221_X1 _18227_ (.A(_06681_),
    .B1(_08937_),
    .B2(_08549_),
    .C1(_08939_),
    .C2(_08631_),
    .ZN(_08940_));
 OAI221_X1 _18228_ (.A(_06695_),
    .B1(_08471_),
    .B2(_08483_),
    .C1(_08736_),
    .C2(_08541_),
    .ZN(_08941_));
 MUX2_X1 _18229_ (.A(_08503_),
    .B(_08468_),
    .S(_08437_),
    .Z(_08942_));
 MUX2_X1 _18230_ (.A(_14792_),
    .B(_08942_),
    .S(_08543_),
    .Z(_08943_));
 OAI21_X1 _18231_ (.A(_08941_),
    .B1(_08943_),
    .B2(_08513_),
    .ZN(_08944_));
 OAI21_X1 _18232_ (.A(_08940_),
    .B1(_08944_),
    .B2(_00396_),
    .ZN(_08945_));
 MUX2_X1 _18233_ (.A(_08935_),
    .B(_08945_),
    .S(_00399_),
    .Z(_08946_));
 NOR2_X1 _18234_ (.A1(net789),
    .A2(_08560_),
    .ZN(_08947_));
 NOR3_X1 _18235_ (.A1(_08483_),
    .A2(_08524_),
    .A3(_08688_),
    .ZN(_08948_));
 OR3_X1 _18236_ (.A1(_08513_),
    .A2(_08947_),
    .A3(_08948_),
    .ZN(_08949_));
 OAI21_X1 _18237_ (.A(_14785_),
    .B1(_08489_),
    .B2(_08493_),
    .ZN(_08950_));
 NAND3_X1 _18238_ (.A1(_00397_),
    .A2(_08615_),
    .A3(_08950_),
    .ZN(_08951_));
 AOI21_X1 _18239_ (.A(_00396_),
    .B1(_08949_),
    .B2(_08951_),
    .ZN(_08952_));
 NOR2_X1 _18240_ (.A1(_14760_),
    .A2(_08560_),
    .ZN(_08953_));
 OAI21_X1 _18241_ (.A(_08536_),
    .B1(_14771_),
    .B2(_14766_),
    .ZN(_08954_));
 OAI22_X1 _18242_ (.A1(_08520_),
    .A2(_00395_),
    .B1(_08953_),
    .B2(_08954_),
    .ZN(_08955_));
 NAND3_X1 _18243_ (.A1(_06681_),
    .A2(_08518_),
    .A3(_08955_),
    .ZN(_08956_));
 OAI21_X1 _18244_ (.A(_08782_),
    .B1(_08915_),
    .B2(_08662_),
    .ZN(_08957_));
 OAI21_X1 _18245_ (.A(_08956_),
    .B1(_08957_),
    .B2(_08518_),
    .ZN(_08958_));
 AOI21_X1 _18246_ (.A(_08736_),
    .B1(_08572_),
    .B2(_08780_),
    .ZN(_08959_));
 OAI21_X1 _18247_ (.A(_08516_),
    .B1(_08914_),
    .B2(_08959_),
    .ZN(_08960_));
 AOI221_X1 _18248_ (.A(_08666_),
    .B1(_08443_),
    .B2(net1124),
    .C1(_08503_),
    .C2(_08499_),
    .ZN(_08961_));
 NAND2_X1 _18249_ (.A1(_08549_),
    .A2(_08961_),
    .ZN(_08962_));
 OAI21_X1 _18250_ (.A(_08478_),
    .B1(_08579_),
    .B2(_08438_),
    .ZN(_08963_));
 OR2_X1 _18251_ (.A1(_08459_),
    .A2(_08963_),
    .ZN(_08964_));
 AND3_X1 _18252_ (.A1(_06681_),
    .A2(_08962_),
    .A3(_08964_),
    .ZN(_08965_));
 OAI22_X1 _18253_ (.A1(_08468_),
    .A2(_08611_),
    .B1(_08799_),
    .B2(_08560_),
    .ZN(_08966_));
 AND3_X1 _18254_ (.A1(_08531_),
    .A2(_08513_),
    .A3(_08966_),
    .ZN(_08967_));
 OAI33_X1 _18255_ (.A1(_08516_),
    .A2(_08952_),
    .A3(_08958_),
    .B1(_08960_),
    .B2(_08965_),
    .B3(_08967_),
    .ZN(_08968_));
 MUX2_X1 _18256_ (.A(_08946_),
    .B(_08968_),
    .S(_00398_),
    .Z(_00031_));
 INV_X1 _18257_ (.A(_06614_),
    .ZN(_08969_));
 BUF_X8 _18258_ (.A(ld_r),
    .Z(_08970_));
 BUF_X16 _18259_ (.A(_08970_),
    .Z(_08971_));
 BUF_X16 _18260_ (.A(_08971_),
    .Z(_08972_));
 BUF_X16 _18261_ (.A(_08972_),
    .Z(_08973_));
 BUF_X16 _18262_ (.A(_08973_),
    .Z(_08974_));
 BUF_X8 _18263_ (.A(_08974_),
    .Z(_08975_));
 NOR2_X2 _18264_ (.A1(_08969_),
    .A2(_08975_),
    .ZN(_08976_));
 NOR2_X2 _18265_ (.A1(_06614_),
    .A2(_08975_),
    .ZN(_08977_));
 BUF_X4 _18266_ (.A(\sa00_sr[7] ),
    .Z(_08978_));
 BUF_X8 _18267_ (.A(\sa10_sr[7] ),
    .Z(_08979_));
 XOR2_X2 _18268_ (.A(_08979_),
    .B(_08978_),
    .Z(_08980_));
 BUF_X4 clone29 (.A(_06351_),
    .Z(net29));
 XOR2_X2 clone8 (.A(_06465_),
    .B(net685),
    .Z(net8));
 XNOR2_X2 _18271_ (.A(\sa20_sr[1] ),
    .B(\sa10_sr[1] ),
    .ZN(_08983_));
 XNOR2_X2 _18272_ (.A(_08983_),
    .B(_08980_),
    .ZN(_08984_));
 BUF_X8 clone36 (.A(net628),
    .Z(net36));
 BUF_X4 _18274_ (.A(\sa10_sr[0] ),
    .Z(_08986_));
 BUF_X8 _18275_ (.A(\sa30_sr[1] ),
    .Z(_08987_));
 XOR2_X2 _18276_ (.A(_08986_),
    .B(_08987_),
    .Z(_08988_));
 XNOR2_X2 _18277_ (.A(\sa00_sr[0] ),
    .B(_08988_),
    .ZN(_08989_));
 XNOR2_X2 _18278_ (.A(_08989_),
    .B(_08984_),
    .ZN(_08990_));
 MUX2_X2 _18279_ (.A(_08976_),
    .B(_08977_),
    .S(_08990_),
    .Z(_08991_));
 BUF_X16 _18280_ (.A(_08970_),
    .Z(_08992_));
 BUF_X8 _18281_ (.A(_08992_),
    .Z(_08993_));
 BUF_X8 _18282_ (.A(_08993_),
    .Z(_08994_));
 BUF_X16 _18283_ (.A(_08994_),
    .Z(_08995_));
 BUF_X8 _18284_ (.A(_08995_),
    .Z(_08996_));
 NOR2_X2 _18285_ (.A1(_06614_),
    .A2(_00440_),
    .ZN(_08997_));
 NAND2_X2 _18286_ (.A1(_08996_),
    .A2(_08997_),
    .ZN(_08998_));
 AND2_X1 _18287_ (.A1(_06614_),
    .A2(_00440_),
    .ZN(_08999_));
 NAND2_X2 _18288_ (.A1(_08996_),
    .A2(_08999_),
    .ZN(_09000_));
 NAND2_X4 _18289_ (.A1(_09000_),
    .A2(_08998_),
    .ZN(_09001_));
 NOR2_X4 _18290_ (.A1(_09001_),
    .A2(_08991_),
    .ZN(_09002_));
 INV_X8 _18291_ (.A(net496),
    .ZN(_09003_));
 BUF_X8 rebuffer421 (.A(_02936_),
    .Z(net884));
 BUF_X16 _18293_ (.A(_09003_),
    .Z(_14800_));
 BUF_X4 clone37 (.A(_09236_),
    .Z(net37));
 BUF_X4 _18295_ (.A(\sa20_sr[0] ),
    .Z(_09006_));
 XNOR2_X2 _18296_ (.A(_08986_),
    .B(_09006_),
    .ZN(_09007_));
 XNOR2_X1 _18297_ (.A(net920),
    .B(_09007_),
    .ZN(_09008_));
 INV_X16 _18298_ (.A(_08970_),
    .ZN(_09009_));
 BUF_X32 _18299_ (.A(_09009_),
    .Z(_09010_));
 BUF_X32 _18300_ (.A(_09010_),
    .Z(_09011_));
 BUF_X32 _18301_ (.A(_09011_),
    .Z(_09012_));
 NAND3_X1 _18302_ (.A1(_06598_),
    .A2(_09012_),
    .A3(net589),
    .ZN(_09013_));
 XNOR2_X2 _18303_ (.A(_08978_),
    .B(_08979_),
    .ZN(_09014_));
 BUF_X16 _18304_ (.A(_08992_),
    .Z(_09015_));
 NOR2_X1 _18305_ (.A1(_06598_),
    .A2(_09015_),
    .ZN(_09016_));
 NAND2_X1 _18306_ (.A1(_09014_),
    .A2(_09016_),
    .ZN(_09017_));
 AOI21_X1 _18307_ (.A(_09008_),
    .B1(_09013_),
    .B2(_09017_),
    .ZN(_09018_));
 XOR2_X2 _18308_ (.A(_08986_),
    .B(_09006_),
    .Z(_09019_));
 XNOR2_X1 _18309_ (.A(net921),
    .B(_09019_),
    .ZN(_09020_));
 NAND2_X1 _18310_ (.A1(net589),
    .A2(_09016_),
    .ZN(_09021_));
 BUF_X8 _18311_ (.A(_09009_),
    .Z(_09022_));
 BUF_X16 _18312_ (.A(_09022_),
    .Z(_09023_));
 NAND3_X1 _18313_ (.A1(_06598_),
    .A2(_09023_),
    .A3(_09014_),
    .ZN(_09024_));
 AOI21_X1 _18314_ (.A(_09020_),
    .B1(_09021_),
    .B2(_09024_),
    .ZN(_09025_));
 INV_X1 _18315_ (.A(_06598_),
    .ZN(_09026_));
 BUF_X16 _18316_ (.A(_08971_),
    .Z(_09027_));
 BUF_X4 _18317_ (.A(_09027_),
    .Z(_09028_));
 NAND3_X1 _18318_ (.A1(_09026_),
    .A2(_09028_),
    .A3(_00441_),
    .ZN(_09029_));
 BUF_X16 _18319_ (.A(_09027_),
    .Z(_09030_));
 NAND2_X1 _18320_ (.A1(_06598_),
    .A2(_09030_),
    .ZN(_09031_));
 OAI21_X1 _18321_ (.A(_09029_),
    .B1(_09031_),
    .B2(_00441_),
    .ZN(_09032_));
 OR3_X4 _18322_ (.A1(_09018_),
    .A2(_09025_),
    .A3(_09032_),
    .ZN(_09033_));
 INV_X4 _18323_ (.A(_09033_),
    .ZN(_09034_));
 BUF_X8 clone561 (.A(net535),
    .Z(net1160));
 BUF_X4 _18325_ (.A(_09034_),
    .Z(_14803_));
 BUF_X8 clone16 (.A(_06225_),
    .Z(net16));
 BUF_X4 _18327_ (.A(\sa30_sr[2] ),
    .Z(_09037_));
 XOR2_X2 _18328_ (.A(\sa10_sr[1] ),
    .B(_09037_),
    .Z(_09038_));
 XOR2_X1 _18329_ (.A(net837),
    .B(_09038_),
    .Z(_09039_));
 BUF_X4 _18330_ (.A(\sa10_sr[2] ),
    .Z(_09040_));
 CLKBUF_X3 _18331_ (.A(\sa20_sr[2] ),
    .Z(_09041_));
 XOR2_X2 _18332_ (.A(_09040_),
    .B(_09041_),
    .Z(_09042_));
 NAND3_X1 _18333_ (.A1(_06630_),
    .A2(_09022_),
    .A3(_09042_),
    .ZN(_09043_));
 XNOR2_X2 _18334_ (.A(_09040_),
    .B(_09041_),
    .ZN(_09044_));
 NOR2_X1 _18335_ (.A1(_06630_),
    .A2(net587),
    .ZN(_09045_));
 NAND2_X1 _18336_ (.A1(_09044_),
    .A2(_09045_),
    .ZN(_09046_));
 AOI21_X2 _18337_ (.A(_09039_),
    .B1(_09043_),
    .B2(_09046_),
    .ZN(_09047_));
 XNOR2_X1 _18338_ (.A(net838),
    .B(_09038_),
    .ZN(_09048_));
 NAND2_X1 _18339_ (.A1(_09042_),
    .A2(_09045_),
    .ZN(_09049_));
 NAND3_X1 _18340_ (.A1(_06630_),
    .A2(net948),
    .A3(_09044_),
    .ZN(_09050_));
 AOI21_X2 _18341_ (.A(_09048_),
    .B1(_09049_),
    .B2(_09050_),
    .ZN(_09051_));
 INV_X1 _18342_ (.A(_06630_),
    .ZN(_09052_));
 NAND3_X1 _18343_ (.A1(_09052_),
    .A2(_08972_),
    .A3(_00442_),
    .ZN(_09053_));
 NAND2_X1 _18344_ (.A1(_06630_),
    .A2(_08972_),
    .ZN(_09054_));
 OAI21_X2 _18345_ (.A(_09053_),
    .B1(_09054_),
    .B2(_00442_),
    .ZN(_09055_));
 NOR3_X4 _18346_ (.A1(_09047_),
    .A2(_09051_),
    .A3(_09055_),
    .ZN(_09056_));
 INV_X4 _18347_ (.A(_09056_),
    .ZN(_09057_));
 BUF_X4 _18348_ (.A(_09057_),
    .Z(_09058_));
 BUF_X4 _18349_ (.A(_09058_),
    .Z(_09059_));
 BUF_X4 _18350_ (.A(_09059_),
    .Z(_09060_));
 BUF_X4 _18351_ (.A(_09060_),
    .Z(_14819_));
 BUF_X8 _18352_ (.A(_09033_),
    .Z(_09061_));
 BUF_X4 _18353_ (.A(_09061_),
    .Z(_14794_));
 BUF_X4 _18354_ (.A(_09056_),
    .Z(_09062_));
 BUF_X4 _18355_ (.A(_09062_),
    .Z(_09063_));
 CLKBUF_X3 _18356_ (.A(_09063_),
    .Z(_09064_));
 BUF_X4 _18357_ (.A(_09064_),
    .Z(_14812_));
 BUF_X2 _18358_ (.A(\sa00_sr[5] ),
    .Z(_09065_));
 BUF_X2 _18359_ (.A(\sa10_sr[6] ),
    .Z(_09066_));
 CLKBUF_X3 _18360_ (.A(\sa20_sr[6] ),
    .Z(_09067_));
 XNOR2_X2 _18361_ (.A(_09066_),
    .B(_09067_),
    .ZN(_09068_));
 XNOR2_X2 _18362_ (.A(_09065_),
    .B(_09068_),
    .ZN(_09069_));
 CLKBUF_X3 _18363_ (.A(\sa10_sr[5] ),
    .Z(_09070_));
 BUF_X4 _18364_ (.A(\sa30_sr[6] ),
    .Z(_09071_));
 XNOR2_X1 _18365_ (.A(_09070_),
    .B(_09071_),
    .ZN(_09072_));
 XNOR2_X1 _18366_ (.A(_09069_),
    .B(_09072_),
    .ZN(_09073_));
 BUF_X8 _18367_ (.A(_09010_),
    .Z(_09074_));
 BUF_X8 _18368_ (.A(_09074_),
    .Z(_09075_));
 BUF_X8 _18369_ (.A(_09075_),
    .Z(_09076_));
 MUX2_X2 _18370_ (.A(\text_in_r[126] ),
    .B(_09073_),
    .S(_09076_),
    .Z(_09077_));
 XOR2_X2 _18371_ (.A(_06701_),
    .B(_09077_),
    .Z(_09078_));
 BUF_X4 _18372_ (.A(_09078_),
    .Z(_09079_));
 BUF_X4 _18373_ (.A(_09079_),
    .Z(_09080_));
 BUF_X4 _18374_ (.A(_09058_),
    .Z(_09081_));
 BUF_X4 _18375_ (.A(_09081_),
    .Z(_09082_));
 BUF_X4 _18376_ (.A(_09082_),
    .Z(_09083_));
 NAND2_X1 _18377_ (.A1(_14794_),
    .A2(_09083_),
    .ZN(_09084_));
 NOR2_X1 _18378_ (.A1(_06649_),
    .A2(_08974_),
    .ZN(_09085_));
 INV_X1 _18379_ (.A(_06649_),
    .ZN(_09086_));
 NOR2_X1 _18380_ (.A1(_09086_),
    .A2(_08974_),
    .ZN(_09087_));
 BUF_X4 _18381_ (.A(\sa00_sr[2] ),
    .Z(_09088_));
 BUF_X2 _18382_ (.A(\sa20_sr[3] ),
    .Z(_09089_));
 XNOR2_X1 _18383_ (.A(_09088_),
    .B(_09089_),
    .ZN(_09090_));
 XNOR2_X2 _18384_ (.A(_08978_),
    .B(_09090_),
    .ZN(_09091_));
 BUF_X2 _18385_ (.A(\sa10_sr[3] ),
    .Z(_09092_));
 XOR2_X2 _18386_ (.A(_08979_),
    .B(_09092_),
    .Z(_09093_));
 BUF_X4 _18387_ (.A(\sa30_sr[3] ),
    .Z(_09094_));
 XNOR2_X1 _18388_ (.A(_09040_),
    .B(_09094_),
    .ZN(_09095_));
 XNOR2_X1 _18389_ (.A(_09093_),
    .B(_09095_),
    .ZN(_09096_));
 XNOR2_X2 _18390_ (.A(_09091_),
    .B(_09096_),
    .ZN(_09097_));
 MUX2_X2 _18391_ (.A(_09085_),
    .B(_09087_),
    .S(_09097_),
    .Z(_09098_));
 BUF_X32 _18392_ (.A(_09010_),
    .Z(_09099_));
 BUF_X16 _18393_ (.A(_09099_),
    .Z(_09100_));
 OR3_X2 _18394_ (.A1(_09086_),
    .A2(net594),
    .A3(\text_in_r[123] ),
    .ZN(_09101_));
 BUF_X16 _18395_ (.A(_09015_),
    .Z(_09102_));
 BUF_X8 _18396_ (.A(_09102_),
    .Z(_09103_));
 NAND3_X2 _18397_ (.A1(_09086_),
    .A2(_09103_),
    .A3(\text_in_r[123] ),
    .ZN(_09104_));
 NAND2_X4 _18398_ (.A1(_09101_),
    .A2(_09104_),
    .ZN(_09105_));
 NOR2_X4 _18399_ (.A1(_09098_),
    .A2(_09105_),
    .ZN(_09106_));
 NOR2_X1 _18400_ (.A1(_09003_),
    .A2(_09106_),
    .ZN(_09107_));
 BUF_X8 _18401_ (.A(_09098_),
    .Z(_09108_));
 OAI21_X4 _18402_ (.A(_09056_),
    .B1(_09108_),
    .B2(_09105_),
    .ZN(_09109_));
 BUF_X4 _18403_ (.A(_14801_),
    .Z(_09110_));
 OAI221_X1 _18404_ (.A(_09080_),
    .B1(_09084_),
    .B2(_09107_),
    .C1(_09109_),
    .C2(_09110_),
    .ZN(_09111_));
 BUF_X4 _18405_ (.A(_09059_),
    .Z(_09112_));
 BUF_X4 _18406_ (.A(_09112_),
    .Z(_09113_));
 CLKBUF_X3 _18407_ (.A(_14804_),
    .Z(_09114_));
 INV_X4 _18408_ (.A(_09114_),
    .ZN(_09115_));
 BUF_X8 _18409_ (.A(_09023_),
    .Z(_09116_));
 NAND2_X1 _18410_ (.A1(_09086_),
    .A2(_09116_),
    .ZN(_09117_));
 BUF_X32 _18411_ (.A(_09012_),
    .Z(_09118_));
 NAND2_X1 _18412_ (.A1(_06649_),
    .A2(_09118_),
    .ZN(_09119_));
 MUX2_X1 _18413_ (.A(_09117_),
    .B(_09119_),
    .S(_09097_),
    .Z(_09120_));
 BUF_X4 _18414_ (.A(_09120_),
    .Z(_09121_));
 BUF_X8 _18415_ (.A(_09121_),
    .Z(_09122_));
 BUF_X4 _18416_ (.A(_09122_),
    .Z(_09123_));
 AND2_X1 _18417_ (.A1(_09101_),
    .A2(_09104_),
    .ZN(_09124_));
 BUF_X4 _18418_ (.A(_09124_),
    .Z(_09125_));
 BUF_X8 _18419_ (.A(_09125_),
    .Z(_09126_));
 BUF_X4 _18420_ (.A(_09126_),
    .Z(_09127_));
 AOI21_X2 _18421_ (.A(_09115_),
    .B1(_09123_),
    .B2(_09127_),
    .ZN(_09128_));
 BUF_X4 _18422_ (.A(_14797_),
    .Z(_09129_));
 BUF_X8 _18423_ (.A(_09105_),
    .Z(_09130_));
 NOR3_X4 _18424_ (.A1(net827),
    .A2(_09108_),
    .A3(_09130_),
    .ZN(_09131_));
 NOR3_X1 _18425_ (.A1(_09113_),
    .A2(_09128_),
    .A3(_09131_),
    .ZN(_09132_));
 BUF_X4 _18426_ (.A(_09106_),
    .Z(_09133_));
 BUF_X4 _18427_ (.A(_09133_),
    .Z(_09134_));
 BUF_X8 _18428_ (.A(_09103_),
    .Z(_09135_));
 BUF_X8 _18429_ (.A(_09135_),
    .Z(_09136_));
 OAI21_X4 _18430_ (.A(_09136_),
    .B1(_08997_),
    .B2(_08999_),
    .ZN(_09137_));
 BUF_X4 _18431_ (.A(_09116_),
    .Z(_09138_));
 NAND2_X1 _18432_ (.A1(_06614_),
    .A2(_09138_),
    .ZN(_09139_));
 NAND2_X1 _18433_ (.A1(_08969_),
    .A2(_09138_),
    .ZN(_09140_));
 MUX2_X2 _18434_ (.A(_09139_),
    .B(_09140_),
    .S(_08990_),
    .Z(_09141_));
 AOI21_X4 _18435_ (.A(_09061_),
    .B1(_09137_),
    .B2(_09141_),
    .ZN(_09142_));
 NAND2_X1 _18436_ (.A1(_09134_),
    .A2(_09142_),
    .ZN(_09143_));
 BUF_X2 split122 (.A(net1147),
    .Z(net122));
 BUF_X4 _18438_ (.A(_09108_),
    .Z(_09145_));
 BUF_X4 _18439_ (.A(_09130_),
    .Z(_09146_));
 OAI21_X2 _18440_ (.A(net1159),
    .B1(_09145_),
    .B2(_09146_),
    .ZN(_09147_));
 AND2_X1 _18441_ (.A1(_09113_),
    .A2(_09147_),
    .ZN(_09148_));
 AOI21_X1 _18442_ (.A(_09132_),
    .B1(_09143_),
    .B2(_09148_),
    .ZN(_09149_));
 OAI21_X1 _18443_ (.A(_09111_),
    .B1(_09149_),
    .B2(_09080_),
    .ZN(_09150_));
 BUF_X8 _18444_ (.A(\sa20_sr[7] ),
    .Z(_09151_));
 BUF_X4 _18445_ (.A(\sa30_sr[7] ),
    .Z(_09152_));
 XOR2_X2 _18446_ (.A(_09152_),
    .B(_09151_),
    .Z(_09153_));
 BUF_X2 _18447_ (.A(\sa00_sr[6] ),
    .Z(_09154_));
 XOR2_X1 _18448_ (.A(_09066_),
    .B(_09154_),
    .Z(_09155_));
 XNOR2_X1 _18449_ (.A(net609),
    .B(_09155_),
    .ZN(_09156_));
 XNOR2_X1 _18450_ (.A(_08979_),
    .B(_09156_),
    .ZN(_09157_));
 BUF_X4 _18451_ (.A(_09076_),
    .Z(_09158_));
 MUX2_X2 _18452_ (.A(\text_in_r[127] ),
    .B(_09157_),
    .S(_09158_),
    .Z(_09159_));
 XNOR2_X2 _18453_ (.A(_06706_),
    .B(_09159_),
    .ZN(_09160_));
 BUF_X2 _18454_ (.A(\sa10_sr[4] ),
    .Z(_09161_));
 BUF_X4 _18455_ (.A(\sa00_sr[4] ),
    .Z(_09162_));
 XNOR2_X2 _18456_ (.A(_09161_),
    .B(_09162_),
    .ZN(_09163_));
 XNOR2_X1 _18457_ (.A(_09070_),
    .B(_09163_),
    .ZN(_09164_));
 BUF_X4 _18458_ (.A(\sa20_sr[5] ),
    .Z(_09165_));
 BUF_X4 _18459_ (.A(\sa30_sr[5] ),
    .Z(_09166_));
 XOR2_X2 _18460_ (.A(_09165_),
    .B(_09166_),
    .Z(_09167_));
 NAND3_X1 _18461_ (.A1(_06683_),
    .A2(_09138_),
    .A3(_09167_),
    .ZN(_09168_));
 XNOR2_X2 _18462_ (.A(_09165_),
    .B(_09166_),
    .ZN(_09169_));
 NOR2_X1 _18463_ (.A1(_06683_),
    .A2(_09103_),
    .ZN(_09170_));
 NAND2_X1 _18464_ (.A1(_09169_),
    .A2(_09170_),
    .ZN(_09171_));
 AOI21_X2 _18465_ (.A(_09164_),
    .B1(_09168_),
    .B2(_09171_),
    .ZN(_09172_));
 XOR2_X1 _18466_ (.A(_09070_),
    .B(_09163_),
    .Z(_09173_));
 NAND2_X1 _18467_ (.A1(_09167_),
    .A2(_09170_),
    .ZN(_09174_));
 BUF_X8 _18468_ (.A(_09116_),
    .Z(_09175_));
 NAND3_X1 _18469_ (.A1(_06683_),
    .A2(_09175_),
    .A3(_09169_),
    .ZN(_09176_));
 AOI21_X2 _18470_ (.A(_09173_),
    .B1(_09174_),
    .B2(_09176_),
    .ZN(_09177_));
 OR3_X1 _18471_ (.A1(_06683_),
    .A2(_09118_),
    .A3(\text_in_r[125] ),
    .ZN(_09178_));
 BUF_X8 _18472_ (.A(_09030_),
    .Z(_09179_));
 BUF_X8 _18473_ (.A(_09179_),
    .Z(_09180_));
 NAND3_X1 _18474_ (.A1(_06683_),
    .A2(_09180_),
    .A3(\text_in_r[125] ),
    .ZN(_09181_));
 NAND2_X1 _18475_ (.A1(_09178_),
    .A2(_09181_),
    .ZN(_09182_));
 NOR3_X4 _18476_ (.A1(_09172_),
    .A2(_09177_),
    .A3(_09182_),
    .ZN(_09183_));
 BUF_X4 _18477_ (.A(_09183_),
    .Z(_09184_));
 CLKBUF_X3 _18478_ (.A(_09184_),
    .Z(_09185_));
 BUF_X2 _18479_ (.A(\sa00_sr[3] ),
    .Z(_09186_));
 BUF_X4 _18480_ (.A(\sa20_sr[4] ),
    .Z(_09187_));
 XNOR2_X1 _18481_ (.A(_09186_),
    .B(_09187_),
    .ZN(_09188_));
 XNOR2_X2 _18482_ (.A(_08978_),
    .B(_09188_),
    .ZN(_09189_));
 BUF_X4 _18483_ (.A(\sa30_sr[4] ),
    .Z(_09190_));
 XOR2_X1 _18484_ (.A(_09161_),
    .B(_09190_),
    .Z(_09191_));
 XNOR2_X1 _18485_ (.A(_09093_),
    .B(_09191_),
    .ZN(_09192_));
 XNOR2_X1 _18486_ (.A(_09189_),
    .B(_09192_),
    .ZN(_09193_));
 BUF_X8 _18487_ (.A(_09022_),
    .Z(_09194_));
 BUF_X8 _18488_ (.A(_09194_),
    .Z(_09195_));
 MUX2_X2 _18489_ (.A(\text_in_r[124] ),
    .B(_09193_),
    .S(_09195_),
    .Z(_09196_));
 XNOR2_X2 _18490_ (.A(_06666_),
    .B(_09196_),
    .ZN(_09197_));
 CLKBUF_X3 _18491_ (.A(_09197_),
    .Z(_09198_));
 CLKBUF_X3 _18492_ (.A(_09198_),
    .Z(_09199_));
 NAND4_X1 _18493_ (.A1(_09150_),
    .A2(_09160_),
    .A3(_09185_),
    .A4(_09199_),
    .ZN(_09200_));
 XNOR2_X2 _18494_ (.A(_06701_),
    .B(_09077_),
    .ZN(_09201_));
 BUF_X4 _18495_ (.A(_09201_),
    .Z(_09202_));
 BUF_X8 _18496_ (.A(_14798_),
    .Z(_09203_));
 NAND3_X2 _18497_ (.A1(_09203_),
    .A2(_09122_),
    .A3(_09126_),
    .ZN(_09204_));
 NAND2_X2 _18498_ (.A1(_09121_),
    .A2(_09125_),
    .ZN(_09205_));
 BUF_X4 _18499_ (.A(_09205_),
    .Z(_09206_));
 BUF_X4 _18500_ (.A(_09206_),
    .Z(_09207_));
 BUF_X4 _18501_ (.A(_09207_),
    .Z(_09208_));
 BUF_X16 _18502_ (.A(_09002_),
    .Z(_09209_));
 BUF_X4 _18503_ (.A(_09209_),
    .Z(_09210_));
 OAI21_X1 _18504_ (.A(_09208_),
    .B1(_14803_),
    .B2(_09210_),
    .ZN(_09211_));
 AOI21_X1 _18505_ (.A(_09083_),
    .B1(_09204_),
    .B2(_09211_),
    .ZN(_09212_));
 XOR2_X2 _18506_ (.A(_06666_),
    .B(_09196_),
    .Z(_09213_));
 BUF_X4 _18507_ (.A(_09213_),
    .Z(_09214_));
 BUF_X4 _18508_ (.A(_09214_),
    .Z(_09215_));
 AOI21_X4 _18509_ (.A(_09062_),
    .B1(_09122_),
    .B2(_09126_),
    .ZN(_09216_));
 CLKBUF_X3 _18510_ (.A(_14806_),
    .Z(_09217_));
 BUF_X8 _18511_ (.A(_09217_),
    .Z(_09218_));
 AOI21_X1 _18512_ (.A(_09215_),
    .B1(_09216_),
    .B2(_09218_),
    .ZN(_09219_));
 INV_X1 _18513_ (.A(_09219_),
    .ZN(_09220_));
 INV_X2 _18514_ (.A(_09203_),
    .ZN(_09221_));
 OAI21_X2 _18515_ (.A(_09214_),
    .B1(_09109_),
    .B2(_09221_),
    .ZN(_09222_));
 NOR2_X4 _18516_ (.A1(_09034_),
    .A2(_09057_),
    .ZN(_09223_));
 AOI221_X1 _18517_ (.A(_09207_),
    .B1(_09223_),
    .B2(_09003_),
    .C1(_09112_),
    .C2(_09114_),
    .ZN(_09224_));
 OAI221_X1 _18518_ (.A(_09202_),
    .B1(_09212_),
    .B2(_09220_),
    .C1(_09222_),
    .C2(_09224_),
    .ZN(_09225_));
 BUF_X4 _18519_ (.A(_09062_),
    .Z(_09226_));
 BUF_X4 _18520_ (.A(_09226_),
    .Z(_09227_));
 AOI21_X2 _18521_ (.A(_09110_),
    .B1(_09123_),
    .B2(_09127_),
    .ZN(_09228_));
 NOR3_X2 _18522_ (.A1(_09203_),
    .A2(_09145_),
    .A3(_09146_),
    .ZN(_09229_));
 OAI21_X1 _18523_ (.A(_09227_),
    .B1(_09228_),
    .B2(_09229_),
    .ZN(_09230_));
 NOR3_X4 _18524_ (.A1(_09062_),
    .A2(_09108_),
    .A3(_09130_),
    .ZN(_09231_));
 NAND2_X1 _18525_ (.A1(net1159),
    .A2(_09231_),
    .ZN(_09232_));
 AND2_X1 _18526_ (.A1(_09230_),
    .A2(_09232_),
    .ZN(_09233_));
 BUF_X4 _18527_ (.A(_09197_),
    .Z(_09234_));
 AOI21_X4 _18528_ (.A(_09081_),
    .B1(_09137_),
    .B2(_09141_),
    .ZN(_09235_));
 INV_X8 _18529_ (.A(_09129_),
    .ZN(_09236_));
 BUF_X16 _18530_ (.A(_09236_),
    .Z(_09237_));
 OAI211_X2 _18531_ (.A(_09123_),
    .B(_09127_),
    .C1(_09237_),
    .C2(_09226_),
    .ZN(_09238_));
 OAI21_X2 _18532_ (.A(_09234_),
    .B1(_09238_),
    .B2(_09235_),
    .ZN(_09239_));
 CLKBUF_X3 _18533_ (.A(_09134_),
    .Z(_09240_));
 NAND2_X4 _18534_ (.A1(_09034_),
    .A2(_09226_),
    .ZN(_09241_));
 NAND2_X1 _18535_ (.A1(_09115_),
    .A2(_09083_),
    .ZN(_09242_));
 AOI21_X1 _18536_ (.A(_09240_),
    .B1(_09241_),
    .B2(_09242_),
    .ZN(_09243_));
 OAI221_X1 _18537_ (.A(_09079_),
    .B1(_09199_),
    .B2(_09233_),
    .C1(_09239_),
    .C2(_09243_),
    .ZN(_09244_));
 AND3_X1 _18538_ (.A1(_09185_),
    .A2(_09225_),
    .A3(_09244_),
    .ZN(_09245_));
 XOR2_X2 _18539_ (.A(_06706_),
    .B(_09159_),
    .Z(_09246_));
 BUF_X4 _18540_ (.A(_09106_),
    .Z(_09247_));
 OAI211_X2 _18541_ (.A(_09061_),
    .B(_09226_),
    .C1(_08991_),
    .C2(_09001_),
    .ZN(_09248_));
 INV_X4 _18542_ (.A(_14801_),
    .ZN(_09249_));
 NAND2_X1 _18543_ (.A1(_09249_),
    .A2(_09058_),
    .ZN(_09250_));
 NAND3_X1 _18544_ (.A1(_09247_),
    .A2(_09248_),
    .A3(_09250_),
    .ZN(_09251_));
 AND2_X1 _18545_ (.A1(_09234_),
    .A2(_09251_),
    .ZN(_09252_));
 OAI21_X4 _18546_ (.A(_09034_),
    .B1(_09108_),
    .B2(_09130_),
    .ZN(_09253_));
 AOI21_X1 _18547_ (.A(_09226_),
    .B1(_09204_),
    .B2(_09253_),
    .ZN(_09254_));
 AOI21_X2 _18548_ (.A(_09057_),
    .B1(_09121_),
    .B2(_09125_),
    .ZN(_09255_));
 BUF_X4 _18549_ (.A(_09255_),
    .Z(_09256_));
 INV_X2 _18550_ (.A(_14796_),
    .ZN(_09257_));
 AOI21_X1 _18551_ (.A(_09254_),
    .B1(_09256_),
    .B2(_09257_),
    .ZN(_09258_));
 BUF_X4 _18552_ (.A(_09247_),
    .Z(_09259_));
 OAI21_X1 _18553_ (.A(_09238_),
    .B1(_09259_),
    .B2(_14817_),
    .ZN(_09260_));
 BUF_X4 _18554_ (.A(_09214_),
    .Z(_09261_));
 AOI221_X1 _18555_ (.A(_09078_),
    .B1(_09252_),
    .B2(_09258_),
    .C1(_09260_),
    .C2(_09261_),
    .ZN(_09262_));
 OR3_X1 _18556_ (.A1(_09172_),
    .A2(_09177_),
    .A3(_09182_),
    .ZN(_09263_));
 BUF_X4 _18557_ (.A(_09263_),
    .Z(_09264_));
 BUF_X4 _18558_ (.A(_09264_),
    .Z(_09265_));
 CLKBUF_X3 _18559_ (.A(_09265_),
    .Z(_09266_));
 CLKBUF_X3 _18560_ (.A(_09266_),
    .Z(_09267_));
 NAND3_X2 _18561_ (.A1(_09217_),
    .A2(_09122_),
    .A3(_09126_),
    .ZN(_09268_));
 OAI21_X4 _18562_ (.A(_09129_),
    .B1(_09108_),
    .B2(_09130_),
    .ZN(_09269_));
 AOI21_X1 _18563_ (.A(_09198_),
    .B1(_09268_),
    .B2(_09269_),
    .ZN(_09270_));
 NOR2_X2 _18564_ (.A1(_09106_),
    .A2(_09213_),
    .ZN(_09271_));
 OAI21_X4 _18565_ (.A(_09034_),
    .B1(_09001_),
    .B2(net525),
    .ZN(_09272_));
 AOI21_X1 _18566_ (.A(_09270_),
    .B1(_09271_),
    .B2(_09272_),
    .ZN(_09273_));
 BUF_X4 _18567_ (.A(_09227_),
    .Z(_09274_));
 NAND2_X1 _18568_ (.A1(_09274_),
    .A2(_09079_),
    .ZN(_09275_));
 NAND2_X1 _18569_ (.A1(_14819_),
    .A2(_09079_),
    .ZN(_09276_));
 AOI21_X4 _18570_ (.A(_09034_),
    .B1(_09121_),
    .B2(_09125_),
    .ZN(_09277_));
 NAND2_X1 _18571_ (.A1(_09234_),
    .A2(_09277_),
    .ZN(_09278_));
 CLKBUF_X3 _18572_ (.A(_09207_),
    .Z(_09279_));
 OAI21_X1 _18573_ (.A(_09278_),
    .B1(_09279_),
    .B2(_09110_),
    .ZN(_09280_));
 OAI221_X1 _18574_ (.A(_09267_),
    .B1(_09273_),
    .B2(_09275_),
    .C1(_09276_),
    .C2(_09280_),
    .ZN(_09281_));
 OAI21_X1 _18575_ (.A(_09246_),
    .B1(_09262_),
    .B2(_09281_),
    .ZN(_09282_));
 NAND3_X2 _18576_ (.A1(_09081_),
    .A2(_09123_),
    .A3(_09127_),
    .ZN(_09283_));
 OAI22_X1 _18577_ (.A1(net37),
    .A2(_09109_),
    .B1(_09283_),
    .B2(_09114_),
    .ZN(_09284_));
 OAI21_X4 _18578_ (.A(_09081_),
    .B1(_09145_),
    .B2(_09146_),
    .ZN(_09285_));
 NAND3_X4 _18579_ (.A1(_09226_),
    .A2(_09123_),
    .A3(_09127_),
    .ZN(_09286_));
 NAND2_X2 _18580_ (.A1(_09285_),
    .A2(_09286_),
    .ZN(_09287_));
 AOI21_X1 _18581_ (.A(_09284_),
    .B1(_09287_),
    .B2(_09257_),
    .ZN(_09288_));
 OAI221_X2 _18582_ (.A(_09079_),
    .B1(_09285_),
    .B2(_14803_),
    .C1(_09286_),
    .C2(_09203_),
    .ZN(_09289_));
 BUF_X2 rebuffer148 (.A(_02272_),
    .Z(net662));
 BUF_X32 _18584_ (.A(_09209_),
    .Z(_14795_));
 AOI21_X1 _18585_ (.A(_09231_),
    .B1(_09256_),
    .B2(_14803_),
    .ZN(_09291_));
 NOR2_X1 _18586_ (.A1(net832),
    .A2(_09291_),
    .ZN(_09292_));
 OAI22_X2 _18587_ (.A1(_09080_),
    .A2(_09288_),
    .B1(_09289_),
    .B2(_09292_),
    .ZN(_09293_));
 NOR2_X2 _18588_ (.A1(_09184_),
    .A2(_09215_),
    .ZN(_09294_));
 NAND3_X4 _18589_ (.A1(_09034_),
    .A2(_09122_),
    .A3(_09126_),
    .ZN(_09295_));
 BUF_X1 split93 (.A(_14810_),
    .Z(net93));
 INV_X2 _18591_ (.A(net826),
    .ZN(_09297_));
 AOI21_X2 _18592_ (.A(_09297_),
    .B1(_09122_),
    .B2(_09126_),
    .ZN(_09298_));
 AOI21_X1 _18593_ (.A(_09298_),
    .B1(_09259_),
    .B2(_09210_),
    .ZN(_09299_));
 OAI221_X1 _18594_ (.A(_09295_),
    .B1(_09109_),
    .B2(net37),
    .C1(_09299_),
    .C2(_09064_),
    .ZN(_09300_));
 NOR2_X4 _18595_ (.A1(_09061_),
    .A2(_09058_),
    .ZN(_09301_));
 AOI21_X1 _18596_ (.A(_09301_),
    .B1(_14794_),
    .B2(_09209_),
    .ZN(_09302_));
 XNOR2_X1 _18597_ (.A(_09259_),
    .B(_09302_),
    .ZN(_09303_));
 MUX2_X1 _18598_ (.A(_09300_),
    .B(_09303_),
    .S(_09202_),
    .Z(_09304_));
 NOR2_X2 _18599_ (.A1(_09264_),
    .A2(_09197_),
    .ZN(_09305_));
 NOR3_X4 _18600_ (.A1(_09237_),
    .A2(_09108_),
    .A3(_09146_),
    .ZN(_09306_));
 NAND2_X1 _18601_ (.A1(_09209_),
    .A2(_09081_),
    .ZN(_09307_));
 NOR2_X2 _18602_ (.A1(_09129_),
    .A2(_09056_),
    .ZN(_09308_));
 NAND2_X1 _18603_ (.A1(_09209_),
    .A2(_09247_),
    .ZN(_09309_));
 AOI221_X2 _18604_ (.A(_09078_),
    .B1(_09306_),
    .B2(_09307_),
    .C1(_09308_),
    .C2(_09309_),
    .ZN(_09310_));
 NOR2_X1 _18605_ (.A1(_09003_),
    .A2(_09208_),
    .ZN(_09311_));
 OAI21_X2 _18606_ (.A(net825),
    .B1(_09145_),
    .B2(_09146_),
    .ZN(_09312_));
 OAI21_X1 _18607_ (.A(_09312_),
    .B1(_09208_),
    .B2(_09210_),
    .ZN(_09313_));
 OAI22_X2 _18608_ (.A1(_09084_),
    .A2(_09311_),
    .B1(_09313_),
    .B2(_09083_),
    .ZN(_09314_));
 AOI21_X1 _18609_ (.A(_09310_),
    .B1(_09314_),
    .B2(_09079_),
    .ZN(_09315_));
 NOR2_X2 _18610_ (.A1(_09184_),
    .A2(_09234_),
    .ZN(_09316_));
 AOI222_X2 _18611_ (.A1(_09293_),
    .A2(_09294_),
    .B1(_09304_),
    .B2(_09305_),
    .C1(_09315_),
    .C2(_09316_),
    .ZN(_09317_));
 OAI221_X2 _18612_ (.A(_09200_),
    .B1(_09245_),
    .B2(_09282_),
    .C1(_09317_),
    .C2(_09246_),
    .ZN(_00032_));
 NOR3_X4 _18613_ (.A1(_09034_),
    .A2(_09098_),
    .A3(_09105_),
    .ZN(_09318_));
 AOI21_X4 _18614_ (.A(_09249_),
    .B1(_09121_),
    .B2(_09125_),
    .ZN(_09319_));
 OAI21_X2 _18615_ (.A(_09064_),
    .B1(_09318_),
    .B2(net870),
    .ZN(_09320_));
 XNOR2_X2 _18616_ (.A(_09003_),
    .B(_09133_),
    .ZN(_09321_));
 OAI211_X2 _18617_ (.A(_09202_),
    .B(_09320_),
    .C1(_09321_),
    .C2(_09274_),
    .ZN(_09322_));
 NOR2_X2 _18618_ (.A1(_09134_),
    .A2(_09272_),
    .ZN(_09323_));
 NAND3_X2 _18619_ (.A1(_09221_),
    .A2(_09123_),
    .A3(_09127_),
    .ZN(_09324_));
 NAND2_X1 _18620_ (.A1(_09082_),
    .A2(_09324_),
    .ZN(_09325_));
 NOR3_X4 _18621_ (.A1(net826),
    .A2(_09098_),
    .A3(_09105_),
    .ZN(_09326_));
 OR2_X4 _18622_ (.A1(_09326_),
    .A2(_09058_),
    .ZN(_09327_));
 AOI21_X4 _18623_ (.A(_09236_),
    .B1(_09121_),
    .B2(_09125_),
    .ZN(_09328_));
 OAI221_X1 _18624_ (.A(_09078_),
    .B1(_09323_),
    .B2(_09325_),
    .C1(_09327_),
    .C2(_09328_),
    .ZN(_09329_));
 AOI21_X1 _18625_ (.A(_09185_),
    .B1(_09329_),
    .B2(_09322_),
    .ZN(_09330_));
 AOI21_X2 _18626_ (.A(_09112_),
    .B1(_09147_),
    .B2(_09324_),
    .ZN(_09331_));
 NOR3_X4 _18627_ (.A1(_09061_),
    .A2(_09108_),
    .A3(_09130_),
    .ZN(_09332_));
 NOR3_X1 _18628_ (.A1(_09227_),
    .A2(_09332_),
    .A3(_09328_),
    .ZN(_09333_));
 NOR3_X1 _18629_ (.A1(_09201_),
    .A2(_09331_),
    .A3(_09333_),
    .ZN(_09334_));
 NOR2_X2 _18630_ (.A1(_09061_),
    .A2(_09062_),
    .ZN(_09335_));
 NOR2_X1 _18631_ (.A1(_09223_),
    .A2(_09335_),
    .ZN(_09336_));
 NOR2_X2 _18632_ (.A1(net497),
    .A2(_09133_),
    .ZN(_09337_));
 NAND2_X1 _18633_ (.A1(net1147),
    .A2(_09081_),
    .ZN(_09338_));
 OAI21_X1 _18634_ (.A(_09338_),
    .B1(_09059_),
    .B2(_09034_),
    .ZN(_09339_));
 AOI221_X2 _18635_ (.A(_09078_),
    .B1(_09336_),
    .B2(_09337_),
    .C1(_09339_),
    .C2(_09134_),
    .ZN(_09340_));
 NOR3_X1 _18636_ (.A1(_09266_),
    .A2(_09334_),
    .A3(_09340_),
    .ZN(_09341_));
 NOR4_X1 _18637_ (.A1(_09341_),
    .A2(_09199_),
    .A3(_09330_),
    .A4(_09246_),
    .ZN(_09342_));
 NOR2_X2 _18638_ (.A1(_09201_),
    .A2(_09265_),
    .ZN(_09343_));
 NOR2_X1 _18639_ (.A1(_09249_),
    .A2(_09081_),
    .ZN(_09344_));
 AOI21_X4 _18640_ (.A(_09062_),
    .B1(_09137_),
    .B2(_09141_),
    .ZN(_09345_));
 OAI21_X1 _18641_ (.A(_09279_),
    .B1(_09344_),
    .B2(_09345_),
    .ZN(_09346_));
 AOI211_X2 _18642_ (.A(_09098_),
    .B(_09130_),
    .C1(_09034_),
    .C2(_09056_),
    .ZN(_09347_));
 NAND2_X1 _18643_ (.A1(_09338_),
    .A2(_09347_),
    .ZN(_09348_));
 NAND3_X1 _18644_ (.A1(_09343_),
    .A2(_09346_),
    .A3(_09348_),
    .ZN(_09349_));
 NAND3_X1 _18645_ (.A1(_09160_),
    .A2(_09199_),
    .A3(_09349_),
    .ZN(_09350_));
 NAND2_X1 _18646_ (.A1(_09078_),
    .A2(_09264_),
    .ZN(_09351_));
 NOR2_X2 _18647_ (.A1(_09206_),
    .A2(_09272_),
    .ZN(_09352_));
 BUF_X16 _18648_ (.A(net827),
    .Z(_09353_));
 AOI21_X2 _18649_ (.A(_09353_),
    .B1(_09123_),
    .B2(_09127_),
    .ZN(_09354_));
 OAI21_X1 _18650_ (.A(_09274_),
    .B1(_09352_),
    .B2(_09354_),
    .ZN(_09355_));
 NAND2_X1 _18651_ (.A1(_14794_),
    .A2(_09231_),
    .ZN(_09356_));
 AOI21_X1 _18652_ (.A(_09351_),
    .B1(_09355_),
    .B2(_09356_),
    .ZN(_09357_));
 NOR2_X1 _18653_ (.A1(_09115_),
    .A2(_09226_),
    .ZN(_09358_));
 NOR2_X1 _18654_ (.A1(_09060_),
    .A2(_09272_),
    .ZN(_09359_));
 NOR3_X1 _18655_ (.A1(_09279_),
    .A2(_09358_),
    .A3(_09359_),
    .ZN(_09360_));
 NOR3_X1 _18656_ (.A1(_14820_),
    .A2(_09240_),
    .A3(_09184_),
    .ZN(_09361_));
 NOR3_X1 _18657_ (.A1(_09079_),
    .A2(_09360_),
    .A3(_09361_),
    .ZN(_09362_));
 NOR2_X1 _18658_ (.A1(_09297_),
    .A2(_09063_),
    .ZN(_09363_));
 NOR2_X1 _18659_ (.A1(_09235_),
    .A2(_09363_),
    .ZN(_09364_));
 NAND2_X1 _18660_ (.A1(_09207_),
    .A2(_09214_),
    .ZN(_09365_));
 NOR3_X4 _18661_ (.A1(_09057_),
    .A2(_09098_),
    .A3(_09105_),
    .ZN(_09366_));
 OAI21_X1 _18662_ (.A(_09366_),
    .B1(_09215_),
    .B2(_09110_),
    .ZN(_09367_));
 OAI221_X1 _18663_ (.A(_09184_),
    .B1(_09364_),
    .B2(_09365_),
    .C1(_09367_),
    .C2(_09142_),
    .ZN(_09368_));
 NOR2_X1 _18664_ (.A1(_09106_),
    .A2(_09142_),
    .ZN(_09369_));
 OAI21_X4 _18665_ (.A(_09237_),
    .B1(_09145_),
    .B2(_09146_),
    .ZN(_09370_));
 NAND3_X1 _18666_ (.A1(_09110_),
    .A2(_09123_),
    .A3(_09127_),
    .ZN(_09371_));
 NAND2_X2 _18667_ (.A1(_09370_),
    .A2(_09371_),
    .ZN(_09372_));
 MUX2_X1 _18668_ (.A(_09369_),
    .B(_09372_),
    .S(_09227_),
    .Z(_09373_));
 AOI21_X2 _18669_ (.A(_09368_),
    .B1(_09373_),
    .B2(_09198_),
    .ZN(_09374_));
 NAND2_X2 _18670_ (.A1(_09078_),
    .A2(_09246_),
    .ZN(_09375_));
 NOR3_X4 _18671_ (.A1(_09257_),
    .A2(_09108_),
    .A3(_09130_),
    .ZN(_09376_));
 NOR3_X2 _18672_ (.A1(_09082_),
    .A2(_09328_),
    .A3(_09376_),
    .ZN(_09377_));
 OAI21_X1 _18673_ (.A(_09112_),
    .B1(_09332_),
    .B2(_09319_),
    .ZN(_09378_));
 NAND2_X1 _18674_ (.A1(_09316_),
    .A2(_09378_),
    .ZN(_09379_));
 OAI22_X1 _18675_ (.A1(_09237_),
    .A2(_09283_),
    .B1(_09253_),
    .B2(_09003_),
    .ZN(_09380_));
 AOI21_X1 _18676_ (.A(_09380_),
    .B1(_09287_),
    .B2(_14794_),
    .ZN(_09381_));
 NAND2_X2 _18677_ (.A1(_09264_),
    .A2(_09197_),
    .ZN(_09382_));
 OAI22_X2 _18678_ (.A1(_09377_),
    .A2(_09379_),
    .B1(_09381_),
    .B2(_09382_),
    .ZN(_09383_));
 OAI33_X1 _18679_ (.A1(_09350_),
    .A2(_09357_),
    .A3(_09362_),
    .B1(_09374_),
    .B2(_09375_),
    .B3(_09383_),
    .ZN(_09384_));
 NAND2_X1 _18680_ (.A1(_09202_),
    .A2(_09246_),
    .ZN(_09385_));
 OAI21_X1 _18681_ (.A(_14800_),
    .B1(_14812_),
    .B2(_09277_),
    .ZN(_09386_));
 NAND2_X4 _18682_ (.A1(_09183_),
    .A2(_09197_),
    .ZN(_09387_));
 AOI221_X1 _18683_ (.A(_09387_),
    .B1(_09318_),
    .B2(net36),
    .C1(_09227_),
    .C2(_09207_),
    .ZN(_09388_));
 OAI21_X4 _18684_ (.A(_09061_),
    .B1(_09108_),
    .B2(_09130_),
    .ZN(_09389_));
 NAND3_X1 _18685_ (.A1(_09083_),
    .A2(_09295_),
    .A3(_09389_),
    .ZN(_09390_));
 AND2_X1 _18686_ (.A1(_09269_),
    .A2(_09371_),
    .ZN(_09391_));
 OAI21_X1 _18687_ (.A(_09390_),
    .B1(_09391_),
    .B2(_09113_),
    .ZN(_09392_));
 AOI22_X1 _18688_ (.A1(_09386_),
    .A2(_09388_),
    .B1(_09392_),
    .B2(_09305_),
    .ZN(_09393_));
 AOI22_X1 _18689_ (.A1(_09249_),
    .A2(_09231_),
    .B1(_09287_),
    .B2(_14800_),
    .ZN(_09394_));
 NAND2_X1 _18690_ (.A1(net831),
    .A2(_09083_),
    .ZN(_09395_));
 NAND2_X1 _18691_ (.A1(net93),
    .A2(_09064_),
    .ZN(_09396_));
 AOI21_X1 _18692_ (.A(_09240_),
    .B1(_09395_),
    .B2(_09396_),
    .ZN(_09397_));
 NAND2_X1 _18693_ (.A1(_09198_),
    .A2(_09251_),
    .ZN(_09398_));
 OAI221_X1 _18694_ (.A(_09267_),
    .B1(_09199_),
    .B2(_09394_),
    .C1(_09397_),
    .C2(_09398_),
    .ZN(_09399_));
 AOI21_X1 _18695_ (.A(_09385_),
    .B1(_09393_),
    .B2(_09399_),
    .ZN(_09400_));
 OR3_X2 _18696_ (.A1(_09384_),
    .A2(_09342_),
    .A3(_09400_),
    .ZN(_00033_));
 NOR2_X1 _18697_ (.A1(_09160_),
    .A2(_09267_),
    .ZN(_09401_));
 NOR2_X1 _18698_ (.A1(_09112_),
    .A2(_09228_),
    .ZN(_09402_));
 AOI21_X4 _18699_ (.A(_09061_),
    .B1(_09121_),
    .B2(_09125_),
    .ZN(_09403_));
 AOI22_X1 _18700_ (.A1(_09114_),
    .A2(_09259_),
    .B1(_09403_),
    .B2(_09003_),
    .ZN(_09404_));
 AOI221_X1 _18701_ (.A(_09222_),
    .B1(_09402_),
    .B2(_09143_),
    .C1(_09404_),
    .C2(_09113_),
    .ZN(_09405_));
 NOR2_X1 _18702_ (.A1(_09354_),
    .A2(_09376_),
    .ZN(_09406_));
 AOI221_X2 _18703_ (.A(_09215_),
    .B1(_09216_),
    .B2(_09110_),
    .C1(_09406_),
    .C2(_09274_),
    .ZN(_09407_));
 NOR3_X1 _18704_ (.A1(_09080_),
    .A2(_09405_),
    .A3(_09407_),
    .ZN(_09408_));
 CLKBUF_X3 _18705_ (.A(_09261_),
    .Z(_09409_));
 NAND2_X1 _18706_ (.A1(_09080_),
    .A2(_09409_),
    .ZN(_09410_));
 NAND3_X1 _18707_ (.A1(net832),
    .A2(_09279_),
    .A3(_09241_),
    .ZN(_09411_));
 NAND2_X1 _18708_ (.A1(_09003_),
    .A2(_09063_),
    .ZN(_09412_));
 MUX2_X1 _18709_ (.A(_09064_),
    .B(_09208_),
    .S(_09003_),
    .Z(_09413_));
 OAI221_X1 _18710_ (.A(_09411_),
    .B1(_09403_),
    .B2(_09412_),
    .C1(net37),
    .C2(_09413_),
    .ZN(_09414_));
 NOR2_X1 _18711_ (.A1(_09240_),
    .A2(_09308_),
    .ZN(_09415_));
 AOI22_X1 _18712_ (.A1(_14817_),
    .A2(_09240_),
    .B1(_09248_),
    .B2(_09415_),
    .ZN(_09416_));
 NAND2_X1 _18713_ (.A1(_09080_),
    .A2(_09199_),
    .ZN(_09417_));
 OAI22_X1 _18714_ (.A1(_09410_),
    .A2(_09414_),
    .B1(_09416_),
    .B2(_09417_),
    .ZN(_09418_));
 OAI21_X1 _18715_ (.A(_09401_),
    .B1(_09408_),
    .B2(_09418_),
    .ZN(_09419_));
 AOI21_X1 _18716_ (.A(_09201_),
    .B1(_14794_),
    .B2(net36),
    .ZN(_09420_));
 INV_X1 _18717_ (.A(_14815_),
    .ZN(_09421_));
 AOI221_X2 _18718_ (.A(_09240_),
    .B1(_09412_),
    .B2(_09420_),
    .C1(_09202_),
    .C2(_09421_),
    .ZN(_09422_));
 NAND2_X1 _18719_ (.A1(_14820_),
    .A2(_09079_),
    .ZN(_09423_));
 NAND4_X1 _18720_ (.A1(_14800_),
    .A2(_14794_),
    .A3(_09113_),
    .A4(_09202_),
    .ZN(_09424_));
 AOI21_X1 _18721_ (.A(_09279_),
    .B1(_09423_),
    .B2(_09424_),
    .ZN(_09425_));
 OAI21_X1 _18722_ (.A(_09199_),
    .B1(_09422_),
    .B2(_09425_),
    .ZN(_09426_));
 NOR3_X1 _18723_ (.A1(_09210_),
    .A2(_09134_),
    .A3(_09335_),
    .ZN(_09427_));
 OAI21_X1 _18724_ (.A(_09202_),
    .B1(_09279_),
    .B2(_14824_),
    .ZN(_09428_));
 NOR3_X1 _18725_ (.A1(_09274_),
    .A2(_09354_),
    .A3(_09376_),
    .ZN(_09429_));
 AOI21_X1 _18726_ (.A(_09128_),
    .B1(_09240_),
    .B2(net832),
    .ZN(_09430_));
 AOI21_X1 _18727_ (.A(_09429_),
    .B1(_09430_),
    .B2(_14812_),
    .ZN(_09431_));
 OAI221_X1 _18728_ (.A(_09409_),
    .B1(_09427_),
    .B2(_09428_),
    .C1(_09431_),
    .C2(_09202_),
    .ZN(_09432_));
 NAND4_X1 _18729_ (.A1(_09246_),
    .A2(_09267_),
    .A3(_09426_),
    .A4(_09432_),
    .ZN(_09433_));
 OAI21_X1 _18730_ (.A(_14819_),
    .B1(_09228_),
    .B2(_09326_),
    .ZN(_09434_));
 NAND3_X1 _18731_ (.A1(_14812_),
    .A2(_09253_),
    .A3(_09268_),
    .ZN(_09435_));
 NAND3_X1 _18732_ (.A1(_09409_),
    .A2(_09434_),
    .A3(_09435_),
    .ZN(_09436_));
 NAND2_X1 _18733_ (.A1(_09274_),
    .A2(_09268_),
    .ZN(_09437_));
 OAI221_X1 _18734_ (.A(_09199_),
    .B1(_09337_),
    .B2(_09437_),
    .C1(_14812_),
    .C2(_09110_),
    .ZN(_09438_));
 NAND4_X1 _18735_ (.A1(_09080_),
    .A2(_09267_),
    .A3(_09436_),
    .A4(_09438_),
    .ZN(_09439_));
 NAND3_X1 _18736_ (.A1(_14812_),
    .A2(_09295_),
    .A3(_09269_),
    .ZN(_09440_));
 NAND3_X1 _18737_ (.A1(_14819_),
    .A2(_09268_),
    .A3(_09370_),
    .ZN(_09441_));
 AOI21_X1 _18738_ (.A(_09409_),
    .B1(_09440_),
    .B2(_09441_),
    .ZN(_09442_));
 NAND3_X2 _18739_ (.A1(net826),
    .A2(_09121_),
    .A3(_09125_),
    .ZN(_09443_));
 OAI211_X2 _18740_ (.A(_14819_),
    .B(_09443_),
    .C1(_09240_),
    .C2(_14800_),
    .ZN(_09444_));
 OAI21_X4 _18741_ (.A(_09218_),
    .B1(_09145_),
    .B2(_09130_),
    .ZN(_09445_));
 NAND3_X1 _18742_ (.A1(_14812_),
    .A2(_09295_),
    .A3(_09445_),
    .ZN(_09446_));
 AOI21_X1 _18743_ (.A(_09199_),
    .B1(_09444_),
    .B2(_09446_),
    .ZN(_09447_));
 OAI21_X1 _18744_ (.A(_09343_),
    .B1(_09442_),
    .B2(_09447_),
    .ZN(_09448_));
 NAND2_X4 _18745_ (.A1(_09183_),
    .A2(_09214_),
    .ZN(_09449_));
 OAI21_X1 _18746_ (.A(_09064_),
    .B1(_09306_),
    .B2(_09403_),
    .ZN(_09450_));
 OAI21_X1 _18747_ (.A(_09221_),
    .B1(_09145_),
    .B2(_09146_),
    .ZN(_09451_));
 OAI211_X2 _18748_ (.A(_09060_),
    .B(_09451_),
    .C1(_09208_),
    .C2(_09210_),
    .ZN(_09452_));
 AOI21_X1 _18749_ (.A(_09449_),
    .B1(_09450_),
    .B2(_09452_),
    .ZN(_09453_));
 NAND2_X4 _18750_ (.A1(_09264_),
    .A2(_09214_),
    .ZN(_09454_));
 NOR3_X2 _18751_ (.A1(_09363_),
    .A2(_09344_),
    .A3(_09207_),
    .ZN(_09455_));
 NOR3_X1 _18752_ (.A1(_09454_),
    .A2(_09427_),
    .A3(_09455_),
    .ZN(_09456_));
 AOI21_X2 _18753_ (.A(_09134_),
    .B1(_09248_),
    .B2(_09250_),
    .ZN(_09457_));
 AND3_X1 _18754_ (.A1(_09295_),
    .A2(_09389_),
    .A3(_09345_),
    .ZN(_09458_));
 NOR2_X1 _18755_ (.A1(net826),
    .A2(_09109_),
    .ZN(_09459_));
 OAI33_X1 _18756_ (.A1(_09239_),
    .A2(_09184_),
    .A3(_09457_),
    .B1(_09458_),
    .B2(_09459_),
    .B3(_09387_),
    .ZN(_09460_));
 OR4_X1 _18757_ (.A1(_09079_),
    .A2(_09460_),
    .A3(_09456_),
    .A4(_09453_),
    .ZN(_09461_));
 NAND4_X1 _18758_ (.A1(_09160_),
    .A2(_09461_),
    .A3(_09448_),
    .A4(_09439_),
    .ZN(_09462_));
 NAND3_X1 _18759_ (.A1(_09419_),
    .A2(_09433_),
    .A3(_09462_),
    .ZN(_00034_));
 NAND3_X1 _18760_ (.A1(_09114_),
    .A2(_09122_),
    .A3(_09126_),
    .ZN(_09463_));
 AOI21_X1 _18761_ (.A(_09059_),
    .B1(_09147_),
    .B2(_09463_),
    .ZN(_09464_));
 NAND3_X2 _18762_ (.A1(_09061_),
    .A2(_09122_),
    .A3(_09126_),
    .ZN(_09465_));
 AOI21_X1 _18763_ (.A(_09063_),
    .B1(_09269_),
    .B2(_09465_),
    .ZN(_09466_));
 AOI211_X2 _18764_ (.A(_09062_),
    .B(_09319_),
    .C1(_09133_),
    .C2(net123),
    .ZN(_09467_));
 NOR3_X1 _18765_ (.A1(_09059_),
    .A2(_09131_),
    .A3(_09298_),
    .ZN(_09468_));
 OAI33_X1 _18766_ (.A1(_09449_),
    .A2(_09464_),
    .A3(_09466_),
    .B1(_09468_),
    .B2(_09467_),
    .B3(_09387_),
    .ZN(_09469_));
 AOI222_X2 _18767_ (.A1(_09353_),
    .A2(_09256_),
    .B1(_09465_),
    .B2(_09345_),
    .C1(_09347_),
    .C2(net124),
    .ZN(_09470_));
 AOI211_X2 _18768_ (.A(_09226_),
    .B(_09328_),
    .C1(_09133_),
    .C2(net123),
    .ZN(_09471_));
 NAND4_X1 _18769_ (.A1(_09061_),
    .A2(_09226_),
    .A3(_09123_),
    .A4(_09127_),
    .ZN(_09472_));
 NAND3_X1 _18770_ (.A1(_09265_),
    .A2(_09214_),
    .A3(_09472_),
    .ZN(_09473_));
 OAI221_X1 _18771_ (.A(_09201_),
    .B1(_09382_),
    .B2(_09470_),
    .C1(_09471_),
    .C2(_09473_),
    .ZN(_09474_));
 OAI21_X1 _18772_ (.A(_09246_),
    .B1(_09469_),
    .B2(_09474_),
    .ZN(_09475_));
 AND3_X1 _18773_ (.A1(_09059_),
    .A2(_09268_),
    .A3(_09312_),
    .ZN(_09476_));
 NAND3_X4 _18774_ (.A1(_09353_),
    .A2(_09122_),
    .A3(_09126_),
    .ZN(_09477_));
 OAI21_X1 _18775_ (.A(_09477_),
    .B1(_09134_),
    .B2(_09003_),
    .ZN(_09478_));
 AOI21_X1 _18776_ (.A(_09476_),
    .B1(_09478_),
    .B2(_09227_),
    .ZN(_09479_));
 NAND2_X2 _18777_ (.A1(_09003_),
    .A2(_09277_),
    .ZN(_09480_));
 AOI21_X1 _18778_ (.A(_09403_),
    .B1(_09247_),
    .B2(_09115_),
    .ZN(_09481_));
 OAI221_X2 _18779_ (.A(_09480_),
    .B1(_09481_),
    .B2(_09063_),
    .C1(net831),
    .C2(_09286_),
    .ZN(_09482_));
 OAI22_X2 _18780_ (.A1(_09454_),
    .A2(_09479_),
    .B1(_09482_),
    .B2(_09449_),
    .ZN(_09483_));
 NAND3_X4 _18781_ (.A1(_09122_),
    .A2(_09126_),
    .A3(_09264_),
    .ZN(_09484_));
 AOI21_X1 _18782_ (.A(_09034_),
    .B1(_09285_),
    .B2(_09484_),
    .ZN(_09485_));
 AOI21_X1 _18783_ (.A(_09485_),
    .B1(_09301_),
    .B2(_09259_),
    .ZN(_09486_));
 AOI22_X2 _18784_ (.A1(_09114_),
    .A2(_09256_),
    .B1(_09231_),
    .B2(net37),
    .ZN(_09487_));
 OAI222_X2 _18785_ (.A1(net832),
    .A2(_09486_),
    .B1(_09487_),
    .B2(_09265_),
    .C1(_09241_),
    .C2(_09484_),
    .ZN(_09488_));
 NOR2_X1 _18786_ (.A1(_09202_),
    .A2(_09261_),
    .ZN(_09489_));
 AOI221_X1 _18787_ (.A(_09475_),
    .B1(_09483_),
    .B2(_09079_),
    .C1(_09488_),
    .C2(_09489_),
    .ZN(_09490_));
 NAND2_X2 _18788_ (.A1(_09078_),
    .A2(_09160_),
    .ZN(_09491_));
 NAND2_X2 _18789_ (.A1(_09221_),
    .A2(_09249_),
    .ZN(_09492_));
 NOR2_X1 _18790_ (.A1(_09247_),
    .A2(_09492_),
    .ZN(_09493_));
 OAI21_X1 _18791_ (.A(_09227_),
    .B1(_09352_),
    .B2(_09493_),
    .ZN(_09494_));
 OAI21_X1 _18792_ (.A(_09463_),
    .B1(_09247_),
    .B2(_09218_),
    .ZN(_09495_));
 AOI21_X1 _18793_ (.A(_09183_),
    .B1(_09495_),
    .B2(_09082_),
    .ZN(_09496_));
 AOI21_X1 _18794_ (.A(_09059_),
    .B1(_09247_),
    .B2(net7),
    .ZN(_09497_));
 OAI222_X2 _18795_ (.A1(net122),
    .A2(_09109_),
    .B1(_09283_),
    .B2(net36),
    .C1(_09497_),
    .C2(_14794_),
    .ZN(_09498_));
 AOI221_X2 _18796_ (.A(_09215_),
    .B1(_09494_),
    .B2(_09496_),
    .C1(_09498_),
    .C2(_09184_),
    .ZN(_09499_));
 NAND2_X4 _18797_ (.A1(_09477_),
    .A2(_09445_),
    .ZN(_09500_));
 OAI221_X1 _18798_ (.A(_09274_),
    .B1(_09265_),
    .B2(_09500_),
    .C1(_09484_),
    .C2(_14803_),
    .ZN(_09501_));
 OAI221_X1 _18799_ (.A(_09083_),
    .B1(_09265_),
    .B2(_09253_),
    .C1(_09279_),
    .C2(net93),
    .ZN(_09502_));
 AND3_X2 _18800_ (.A1(_09409_),
    .A2(_09501_),
    .A3(_09502_),
    .ZN(_09503_));
 NAND2_X2 _18801_ (.A1(_09202_),
    .A2(_09160_),
    .ZN(_09504_));
 NOR2_X1 _18802_ (.A1(_09216_),
    .A2(_09366_),
    .ZN(_09505_));
 AOI221_X2 _18803_ (.A(_09387_),
    .B1(_09301_),
    .B2(_09259_),
    .C1(_09505_),
    .C2(_09218_),
    .ZN(_09506_));
 NOR3_X1 _18804_ (.A1(_09113_),
    .A2(_09131_),
    .A3(_09493_),
    .ZN(_09507_));
 OAI21_X1 _18805_ (.A(_09059_),
    .B1(_09332_),
    .B2(_09298_),
    .ZN(_09508_));
 NAND2_X1 _18806_ (.A1(_09294_),
    .A2(_09508_),
    .ZN(_09509_));
 OR3_X1 _18807_ (.A1(_09235_),
    .A2(_09358_),
    .A3(_09484_),
    .ZN(_09510_));
 NOR4_X1 _18808_ (.A1(_09059_),
    .A2(_09145_),
    .A3(_09146_),
    .A4(_09264_),
    .ZN(_09511_));
 NOR2_X1 _18809_ (.A1(_09063_),
    .A2(_09184_),
    .ZN(_09512_));
 AOI21_X1 _18810_ (.A(_09511_),
    .B1(_09512_),
    .B2(_09207_),
    .ZN(_09513_));
 OAI21_X1 _18811_ (.A(_09510_),
    .B1(_09513_),
    .B2(net831),
    .ZN(_09514_));
 OAI22_X1 _18812_ (.A1(_09507_),
    .A2(_09509_),
    .B1(_09514_),
    .B2(_09222_),
    .ZN(_09515_));
 OAI33_X1 _18813_ (.A1(_09503_),
    .A2(_09499_),
    .A3(_09491_),
    .B1(_09504_),
    .B2(_09506_),
    .B3(_09515_),
    .ZN(_09516_));
 OR2_X1 _18814_ (.A1(_09516_),
    .A2(_09490_),
    .ZN(_00035_));
 AOI22_X1 _18815_ (.A1(_09297_),
    .A2(_09231_),
    .B1(_09465_),
    .B2(_09274_),
    .ZN(_09517_));
 NOR2_X1 _18816_ (.A1(_09382_),
    .A2(_09517_),
    .ZN(_09518_));
 NOR2_X1 _18817_ (.A1(_09229_),
    .A2(_09323_),
    .ZN(_09519_));
 NOR3_X1 _18818_ (.A1(_14812_),
    .A2(_09449_),
    .A3(_09519_),
    .ZN(_09520_));
 NOR2_X1 _18819_ (.A1(_09110_),
    .A2(_09207_),
    .ZN(_09521_));
 NOR3_X1 _18820_ (.A1(_09060_),
    .A2(_09521_),
    .A3(_09323_),
    .ZN(_09522_));
 NOR3_X2 _18821_ (.A1(_09064_),
    .A2(_09306_),
    .A3(_09277_),
    .ZN(_09523_));
 NOR3_X1 _18822_ (.A1(_09060_),
    .A2(_09228_),
    .A3(_09376_),
    .ZN(_09524_));
 NOR2_X1 _18823_ (.A1(_09227_),
    .A2(_09321_),
    .ZN(_09525_));
 OAI33_X1 _18824_ (.A1(_09523_),
    .A2(_09522_),
    .A3(_09387_),
    .B1(_09524_),
    .B2(_09525_),
    .B3(_09454_),
    .ZN(_09526_));
 OR4_X2 _18825_ (.A1(_09526_),
    .A2(_09518_),
    .A3(_09520_),
    .A4(_09491_),
    .ZN(_09527_));
 NAND2_X1 _18826_ (.A1(_09082_),
    .A2(_09445_),
    .ZN(_09528_));
 NAND2_X1 _18827_ (.A1(net123),
    .A2(_09318_),
    .ZN(_09529_));
 NAND2_X1 _18828_ (.A1(net832),
    .A2(_09256_),
    .ZN(_09530_));
 NAND4_X1 _18829_ (.A1(_09305_),
    .A2(_09528_),
    .A3(_09529_),
    .A4(_09530_),
    .ZN(_09531_));
 OAI21_X1 _18830_ (.A(_09060_),
    .B1(_09403_),
    .B2(_09376_),
    .ZN(_09532_));
 OAI221_X2 _18831_ (.A(_09532_),
    .B1(_09389_),
    .B2(net832),
    .C1(_09203_),
    .C2(_09286_),
    .ZN(_09533_));
 NOR2_X1 _18832_ (.A1(_14808_),
    .A2(_09208_),
    .ZN(_09534_));
 AOI21_X2 _18833_ (.A(_09534_),
    .B1(_09395_),
    .B2(_09279_),
    .ZN(_09535_));
 OAI221_X2 _18834_ (.A(_09531_),
    .B1(_09533_),
    .B2(_09382_),
    .C1(_09387_),
    .C2(_09535_),
    .ZN(_09536_));
 INV_X2 _18835_ (.A(_09217_),
    .ZN(_09537_));
 NOR2_X1 _18836_ (.A1(_09277_),
    .A2(_09311_),
    .ZN(_09538_));
 OAI221_X1 _18837_ (.A(_09143_),
    .B1(_09285_),
    .B2(_09537_),
    .C1(_09538_),
    .C2(_14819_),
    .ZN(_09539_));
 AOI21_X1 _18838_ (.A(_09536_),
    .B1(_09539_),
    .B2(_09316_),
    .ZN(_09540_));
 AND2_X1 _18839_ (.A1(_14819_),
    .A2(_09391_),
    .ZN(_09541_));
 OAI21_X1 _18840_ (.A(_09185_),
    .B1(_14819_),
    .B2(_09218_),
    .ZN(_09542_));
 AOI221_X1 _18841_ (.A(_09082_),
    .B1(_09134_),
    .B2(_09249_),
    .C1(_09277_),
    .C2(_09003_),
    .ZN(_09543_));
 AOI21_X2 _18842_ (.A(_09326_),
    .B1(_09206_),
    .B2(net7),
    .ZN(_09544_));
 AOI21_X1 _18843_ (.A(_09543_),
    .B1(_09544_),
    .B2(_14819_),
    .ZN(_09545_));
 OAI221_X1 _18844_ (.A(_09409_),
    .B1(_09541_),
    .B2(_09542_),
    .C1(_09545_),
    .C2(_09185_),
    .ZN(_09546_));
 NOR2_X1 _18845_ (.A1(_09112_),
    .A2(_09326_),
    .ZN(_09547_));
 AOI221_X2 _18846_ (.A(_09387_),
    .B1(_09547_),
    .B2(_09480_),
    .C1(_09500_),
    .C2(_09083_),
    .ZN(_09548_));
 NOR2_X1 _18847_ (.A1(net122),
    .A2(_09112_),
    .ZN(_09549_));
 OAI21_X1 _18848_ (.A(_09208_),
    .B1(_09345_),
    .B2(_09549_),
    .ZN(_09550_));
 AND4_X1 _18849_ (.A1(_09266_),
    .A2(_09198_),
    .A3(_09251_),
    .A4(_09550_),
    .ZN(_09551_));
 NOR2_X1 _18850_ (.A1(_09548_),
    .A2(_09551_),
    .ZN(_09552_));
 AOI21_X1 _18851_ (.A(_09080_),
    .B1(_09546_),
    .B2(_09552_),
    .ZN(_09553_));
 NAND2_X1 _18852_ (.A1(_09324_),
    .A2(_09528_),
    .ZN(_09554_));
 OR3_X1 _18853_ (.A1(_09227_),
    .A2(_09337_),
    .A3(_09376_),
    .ZN(_09555_));
 NOR2_X1 _18854_ (.A1(_09261_),
    .A2(_09301_),
    .ZN(_09556_));
 AOI221_X2 _18855_ (.A(_09266_),
    .B1(_09261_),
    .B2(_09554_),
    .C1(_09555_),
    .C2(_09556_),
    .ZN(_09557_));
 NOR2_X1 _18856_ (.A1(net832),
    .A2(_09287_),
    .ZN(_09558_));
 OAI221_X2 _18857_ (.A(_09294_),
    .B1(_09241_),
    .B2(_09208_),
    .C1(_14800_),
    .C2(_09389_),
    .ZN(_09559_));
 OAI221_X2 _18858_ (.A(_09316_),
    .B1(_09113_),
    .B2(_14800_),
    .C1(_09257_),
    .C2(_09285_),
    .ZN(_09560_));
 OAI221_X2 _18859_ (.A(_09080_),
    .B1(_09558_),
    .B2(_09559_),
    .C1(_09560_),
    .C2(_09352_),
    .ZN(_09561_));
 OAI21_X1 _18860_ (.A(_09246_),
    .B1(_09557_),
    .B2(_09561_),
    .ZN(_09562_));
 OAI221_X1 _18861_ (.A(_09527_),
    .B1(_09540_),
    .B2(_09504_),
    .C1(_09553_),
    .C2(_09562_),
    .ZN(_00036_));
 NAND2_X1 _18862_ (.A1(_09204_),
    .A2(_09269_),
    .ZN(_09563_));
 AOI221_X2 _18863_ (.A(_09234_),
    .B1(_09366_),
    .B2(net36),
    .C1(_09563_),
    .C2(_09060_),
    .ZN(_09564_));
 OAI21_X1 _18864_ (.A(_09443_),
    .B1(_09247_),
    .B2(net1159),
    .ZN(_09565_));
 AOI221_X1 _18865_ (.A(_09215_),
    .B1(_09565_),
    .B2(_09082_),
    .C1(_09256_),
    .C2(net37),
    .ZN(_09566_));
 NOR3_X1 _18866_ (.A1(_09185_),
    .A2(_09564_),
    .A3(_09566_),
    .ZN(_09567_));
 AOI22_X1 _18867_ (.A1(_09114_),
    .A2(_09216_),
    .B1(_09366_),
    .B2(_14794_),
    .ZN(_09568_));
 NAND2_X1 _18868_ (.A1(_14795_),
    .A2(_09198_),
    .ZN(_09569_));
 OAI221_X1 _18869_ (.A(_09185_),
    .B1(_09198_),
    .B2(_09568_),
    .C1(_09569_),
    .C2(_09231_),
    .ZN(_09570_));
 NOR2_X1 _18870_ (.A1(_09256_),
    .A2(_09198_),
    .ZN(_09571_));
 NAND2_X1 _18871_ (.A1(net628),
    .A2(_09214_),
    .ZN(_09572_));
 OAI33_X1 _18872_ (.A1(net832),
    .A2(_09271_),
    .A3(_09571_),
    .B1(_09572_),
    .B2(_09146_),
    .B3(_09145_),
    .ZN(_09573_));
 AOI21_X1 _18873_ (.A(_09570_),
    .B1(_09573_),
    .B2(_14803_),
    .ZN(_09574_));
 NOR4_X1 _18874_ (.A1(_09210_),
    .A2(_09207_),
    .A3(_09223_),
    .A4(_09335_),
    .ZN(_09575_));
 NOR2_X1 _18875_ (.A1(_09203_),
    .A2(_09110_),
    .ZN(_09576_));
 OAI21_X1 _18876_ (.A(_09576_),
    .B1(_09146_),
    .B2(_09145_),
    .ZN(_09577_));
 NOR2_X1 _18877_ (.A1(_09060_),
    .A2(_09577_),
    .ZN(_09578_));
 OR3_X1 _18878_ (.A1(_09261_),
    .A2(_09575_),
    .A3(_09578_),
    .ZN(_09579_));
 NOR2_X1 _18879_ (.A1(_09249_),
    .A2(_09064_),
    .ZN(_09580_));
 OAI221_X1 _18880_ (.A(_09261_),
    .B1(_09285_),
    .B2(net93),
    .C1(_09580_),
    .C2(_09279_),
    .ZN(_09581_));
 AOI21_X1 _18881_ (.A(_09267_),
    .B1(_09579_),
    .B2(_09581_),
    .ZN(_09582_));
 AOI21_X1 _18882_ (.A(_09128_),
    .B1(_09142_),
    .B2(_09366_),
    .ZN(_09583_));
 OAI21_X1 _18883_ (.A(_09266_),
    .B1(_09261_),
    .B2(_09583_),
    .ZN(_09584_));
 NOR3_X1 _18884_ (.A1(_09083_),
    .A2(_09306_),
    .A3(_09354_),
    .ZN(_09585_));
 NOR2_X1 _18885_ (.A1(_09128_),
    .A2(_09326_),
    .ZN(_09586_));
 AOI21_X1 _18886_ (.A(_09585_),
    .B1(_09586_),
    .B2(_09113_),
    .ZN(_09587_));
 AOI21_X1 _18887_ (.A(_09584_),
    .B1(_09587_),
    .B2(_09409_),
    .ZN(_09588_));
 OAI33_X1 _18888_ (.A1(_09385_),
    .A2(_09567_),
    .A3(_09574_),
    .B1(_09588_),
    .B2(_09582_),
    .B3(_09504_),
    .ZN(_09589_));
 NOR2_X1 _18889_ (.A1(_14819_),
    .A2(_09500_),
    .ZN(_09590_));
 OAI21_X1 _18890_ (.A(_09266_),
    .B1(_09253_),
    .B2(_09274_),
    .ZN(_09591_));
 OAI21_X1 _18891_ (.A(_09312_),
    .B1(_09279_),
    .B2(_14800_),
    .ZN(_09592_));
 OAI21_X1 _18892_ (.A(_09230_),
    .B1(_09592_),
    .B2(_14812_),
    .ZN(_09593_));
 OAI221_X1 _18893_ (.A(_09199_),
    .B1(_09590_),
    .B2(_09591_),
    .C1(_09593_),
    .C2(_09267_),
    .ZN(_09594_));
 AOI221_X2 _18894_ (.A(_09206_),
    .B1(_09223_),
    .B2(_09003_),
    .C1(_09082_),
    .C2(_09537_),
    .ZN(_09595_));
 NOR4_X1 _18895_ (.A1(_09267_),
    .A2(_09222_),
    .A3(net871),
    .A4(_09595_),
    .ZN(_09596_));
 NAND2_X1 _18896_ (.A1(_14812_),
    .A2(_09371_),
    .ZN(_09597_));
 AOI21_X1 _18897_ (.A(_09454_),
    .B1(_09480_),
    .B2(_09597_),
    .ZN(_09598_));
 NOR2_X1 _18898_ (.A1(_09596_),
    .A2(_09598_),
    .ZN(_09599_));
 AOI21_X1 _18899_ (.A(_09375_),
    .B1(_09594_),
    .B2(_09599_),
    .ZN(_09600_));
 NOR2_X1 _18900_ (.A1(net628),
    .A2(_09206_),
    .ZN(_09601_));
 NOR3_X1 _18901_ (.A1(_14803_),
    .A2(_09265_),
    .A3(_09601_),
    .ZN(_09602_));
 NOR2_X1 _18902_ (.A1(_09261_),
    .A2(_09602_),
    .ZN(_09603_));
 OAI221_X1 _18903_ (.A(_09112_),
    .B1(_09259_),
    .B2(_09034_),
    .C1(_09484_),
    .C2(_09110_),
    .ZN(_09604_));
 NAND4_X1 _18904_ (.A1(_09003_),
    .A2(_09034_),
    .A3(_09206_),
    .A4(_09265_),
    .ZN(_09605_));
 NAND2_X1 _18905_ (.A1(_09034_),
    .A2(_09183_),
    .ZN(_09606_));
 OAI221_X1 _18906_ (.A(_09605_),
    .B1(_09606_),
    .B2(_09207_),
    .C1(_09484_),
    .C2(_14803_),
    .ZN(_09607_));
 OAI21_X1 _18907_ (.A(_09604_),
    .B1(_09607_),
    .B2(_09083_),
    .ZN(_09608_));
 AOI21_X1 _18908_ (.A(_09062_),
    .B1(_09133_),
    .B2(_09537_),
    .ZN(_09609_));
 OAI21_X1 _18909_ (.A(_09269_),
    .B1(_09206_),
    .B2(net7),
    .ZN(_09610_));
 AOI221_X2 _18910_ (.A(_09264_),
    .B1(_09480_),
    .B2(_09609_),
    .C1(_09610_),
    .C2(_09063_),
    .ZN(_09611_));
 AOI22_X1 _18911_ (.A1(_09272_),
    .A2(_09366_),
    .B1(_09586_),
    .B2(_09060_),
    .ZN(_09612_));
 AOI21_X1 _18912_ (.A(_09611_),
    .B1(_09612_),
    .B2(_09266_),
    .ZN(_09613_));
 AOI221_X2 _18913_ (.A(_09491_),
    .B1(_09603_),
    .B2(_09608_),
    .C1(_09613_),
    .C2(_09409_),
    .ZN(_09614_));
 NOR3_X1 _18914_ (.A1(_09589_),
    .A2(_09600_),
    .A3(_09614_),
    .ZN(_00037_));
 INV_X1 _18915_ (.A(_09504_),
    .ZN(_09615_));
 NOR2_X1 _18916_ (.A1(_09409_),
    .A2(_09457_),
    .ZN(_09616_));
 AOI221_X2 _18917_ (.A(_09198_),
    .B1(_09495_),
    .B2(_09082_),
    .C1(_09256_),
    .C2(_09210_),
    .ZN(_09617_));
 NOR3_X1 _18918_ (.A1(_09185_),
    .A2(_09616_),
    .A3(_09617_),
    .ZN(_09618_));
 OAI21_X1 _18919_ (.A(_09508_),
    .B1(_09109_),
    .B2(net831),
    .ZN(_09619_));
 AOI21_X1 _18920_ (.A(_09215_),
    .B1(_09208_),
    .B2(_14814_),
    .ZN(_09620_));
 NAND2_X1 _18921_ (.A1(_09218_),
    .A2(_09112_),
    .ZN(_09621_));
 NAND3_X1 _18922_ (.A1(_09259_),
    .A2(_09412_),
    .A3(_09621_),
    .ZN(_09622_));
 AOI221_X2 _18923_ (.A(_09265_),
    .B1(_09261_),
    .B2(_09619_),
    .C1(_09620_),
    .C2(_09622_),
    .ZN(_09623_));
 OAI21_X1 _18924_ (.A(_09615_),
    .B1(_09618_),
    .B2(_09623_),
    .ZN(_09624_));
 AOI21_X1 _18925_ (.A(_09335_),
    .B1(_09277_),
    .B2(net628),
    .ZN(_09625_));
 AOI21_X1 _18926_ (.A(_09332_),
    .B1(_09223_),
    .B2(net628),
    .ZN(_09626_));
 OAI21_X1 _18927_ (.A(_09625_),
    .B1(_09626_),
    .B2(net93),
    .ZN(_09627_));
 OAI21_X1 _18928_ (.A(_09063_),
    .B1(_09234_),
    .B2(_09326_),
    .ZN(_09628_));
 OAI21_X1 _18929_ (.A(_09628_),
    .B1(_09215_),
    .B2(_14803_),
    .ZN(_09629_));
 AOI222_X2 _18930_ (.A1(_09301_),
    .A2(_09271_),
    .B1(_09627_),
    .B2(_09215_),
    .C1(_14800_),
    .C2(_09629_),
    .ZN(_09630_));
 OR3_X1 _18931_ (.A1(_09267_),
    .A2(_09491_),
    .A3(_09630_),
    .ZN(_09631_));
 NAND2_X4 _18932_ (.A1(_09353_),
    .A2(_09197_),
    .ZN(_09632_));
 AOI221_X2 _18933_ (.A(_09081_),
    .B1(_09133_),
    .B2(_09632_),
    .C1(_09271_),
    .C2(_09537_),
    .ZN(_09633_));
 AOI21_X1 _18934_ (.A(_09227_),
    .B1(_09278_),
    .B2(_09572_),
    .ZN(_09634_));
 NOR3_X1 _18935_ (.A1(_09201_),
    .A2(_09246_),
    .A3(_09183_),
    .ZN(_09635_));
 OAI21_X1 _18936_ (.A(_09635_),
    .B1(_09234_),
    .B2(_09295_),
    .ZN(_09636_));
 NOR3_X2 _18937_ (.A1(_09634_),
    .A2(_09633_),
    .A3(_09636_),
    .ZN(_09637_));
 NOR2_X1 _18938_ (.A1(_09184_),
    .A2(_09375_),
    .ZN(_09638_));
 AOI21_X1 _18939_ (.A(_09057_),
    .B1(_09205_),
    .B2(_09203_),
    .ZN(_09639_));
 OAI22_X2 _18940_ (.A1(_09217_),
    .A2(_09205_),
    .B1(_09253_),
    .B2(net496),
    .ZN(_09640_));
 AOI221_X2 _18941_ (.A(_09213_),
    .B1(_09443_),
    .B2(_09639_),
    .C1(_09640_),
    .C2(_09058_),
    .ZN(_09641_));
 NAND3_X1 _18942_ (.A1(_09059_),
    .A2(_09477_),
    .A3(_09577_),
    .ZN(_09642_));
 OAI21_X1 _18943_ (.A(_09295_),
    .B1(_09134_),
    .B2(_09218_),
    .ZN(_09643_));
 OAI21_X1 _18944_ (.A(_09642_),
    .B1(_09643_),
    .B2(_09082_),
    .ZN(_09644_));
 AOI21_X1 _18945_ (.A(_09641_),
    .B1(_09644_),
    .B2(_09215_),
    .ZN(_09645_));
 NAND2_X1 _18946_ (.A1(net496),
    .A2(_09062_),
    .ZN(_09646_));
 NOR2_X1 _18947_ (.A1(_14813_),
    .A2(_14822_),
    .ZN(_09647_));
 AOI221_X1 _18948_ (.A(_09213_),
    .B1(_09369_),
    .B2(_09646_),
    .C1(_09647_),
    .C2(_09133_),
    .ZN(_09648_));
 NOR3_X1 _18949_ (.A1(_09266_),
    .A2(_09375_),
    .A3(_09648_),
    .ZN(_09649_));
 OAI21_X1 _18950_ (.A(_09445_),
    .B1(_09206_),
    .B2(net122),
    .ZN(_09650_));
 AOI22_X1 _18951_ (.A1(_09203_),
    .A2(_09216_),
    .B1(_09650_),
    .B2(_09063_),
    .ZN(_09651_));
 OR2_X1 _18952_ (.A1(_09198_),
    .A2(_09651_),
    .ZN(_09652_));
 AOI221_X2 _18953_ (.A(_09637_),
    .B1(_09638_),
    .B2(_09645_),
    .C1(_09649_),
    .C2(_09652_),
    .ZN(_09653_));
 NOR3_X1 _18954_ (.A1(_09210_),
    .A2(_14803_),
    .A3(_09064_),
    .ZN(_09654_));
 OAI21_X1 _18955_ (.A(_09259_),
    .B1(_09060_),
    .B2(_09353_),
    .ZN(_09655_));
 NOR3_X1 _18956_ (.A1(_09449_),
    .A2(_09654_),
    .A3(_09655_),
    .ZN(_09656_));
 NOR3_X1 _18957_ (.A1(_14815_),
    .A2(_09240_),
    .A3(_09449_),
    .ZN(_09657_));
 NOR3_X1 _18958_ (.A1(_09385_),
    .A2(_09656_),
    .A3(_09657_),
    .ZN(_09658_));
 AOI21_X1 _18959_ (.A(_09240_),
    .B1(_09241_),
    .B2(_14800_),
    .ZN(_09659_));
 AOI21_X1 _18960_ (.A(_09659_),
    .B1(_09231_),
    .B2(_09115_),
    .ZN(_09660_));
 NOR2_X1 _18961_ (.A1(_09210_),
    .A2(_09389_),
    .ZN(_09661_));
 OAI21_X1 _18962_ (.A(_09064_),
    .B1(_09208_),
    .B2(_09492_),
    .ZN(_09662_));
 NAND2_X1 _18963_ (.A1(_09477_),
    .A2(_09253_),
    .ZN(_09663_));
 OAI221_X1 _18964_ (.A(_09266_),
    .B1(_09661_),
    .B2(_09662_),
    .C1(_09663_),
    .C2(_09274_),
    .ZN(_09664_));
 OAI22_X1 _18965_ (.A1(_09113_),
    .A2(_09478_),
    .B1(_09661_),
    .B2(_09325_),
    .ZN(_09665_));
 OAI21_X1 _18966_ (.A(_09664_),
    .B1(_09665_),
    .B2(_09267_),
    .ZN(_09666_));
 OAI221_X1 _18967_ (.A(_09658_),
    .B1(_09660_),
    .B2(_09454_),
    .C1(_09409_),
    .C2(_09666_),
    .ZN(_09667_));
 AND4_X2 _18968_ (.A1(_09631_),
    .A2(_09653_),
    .A3(_09624_),
    .A4(_09667_),
    .ZN(_00038_));
 AOI21_X1 _18969_ (.A(_09459_),
    .B1(_09318_),
    .B2(_09081_),
    .ZN(_09668_));
 AOI221_X2 _18970_ (.A(_09197_),
    .B1(_09366_),
    .B2(_09236_),
    .C1(_09308_),
    .C2(_09205_),
    .ZN(_09669_));
 OAI21_X1 _18971_ (.A(_09058_),
    .B1(_09206_),
    .B2(_09218_),
    .ZN(_09670_));
 OAI22_X2 _18972_ (.A1(_09277_),
    .A2(_09327_),
    .B1(_09670_),
    .B2(_09107_),
    .ZN(_09671_));
 AOI221_X2 _18973_ (.A(_09351_),
    .B1(_09668_),
    .B2(_09669_),
    .C1(_09671_),
    .C2(_09234_),
    .ZN(_09672_));
 NOR4_X1 _18974_ (.A1(net7),
    .A2(_09034_),
    .A3(_09109_),
    .A4(_09197_),
    .ZN(_09673_));
 OAI21_X1 _18975_ (.A(_09283_),
    .B1(_09214_),
    .B2(_09134_),
    .ZN(_09674_));
 AOI21_X1 _18976_ (.A(_09673_),
    .B1(_09674_),
    .B2(_09142_),
    .ZN(_09675_));
 AOI221_X1 _18977_ (.A(_09183_),
    .B1(_09197_),
    .B2(_09058_),
    .C1(_09366_),
    .C2(net831),
    .ZN(_09676_));
 AOI21_X1 _18978_ (.A(_09078_),
    .B1(_09675_),
    .B2(_09676_),
    .ZN(_09677_));
 OAI21_X1 _18979_ (.A(net7),
    .B1(_09231_),
    .B2(_09403_),
    .ZN(_09678_));
 AOI21_X1 _18980_ (.A(_09214_),
    .B1(_09529_),
    .B2(_09678_),
    .ZN(_09679_));
 AOI21_X1 _18981_ (.A(_09332_),
    .B1(_09256_),
    .B2(_14794_),
    .ZN(_09680_));
 AOI21_X1 _18982_ (.A(_09216_),
    .B1(_09301_),
    .B2(_09247_),
    .ZN(_09681_));
 OAI22_X1 _18983_ (.A1(_09234_),
    .A2(_09680_),
    .B1(_09681_),
    .B2(net36),
    .ZN(_09682_));
 OAI21_X1 _18984_ (.A(_09184_),
    .B1(_09679_),
    .B2(_09682_),
    .ZN(_09683_));
 OAI221_X1 _18985_ (.A(_09234_),
    .B1(_09285_),
    .B2(_09218_),
    .C1(_09544_),
    .C2(_09112_),
    .ZN(_09684_));
 AOI221_X2 _18986_ (.A(_09197_),
    .B1(_09318_),
    .B2(_09058_),
    .C1(_09255_),
    .C2(net122),
    .ZN(_09685_));
 OAI221_X1 _18987_ (.A(_09685_),
    .B1(_09285_),
    .B2(_09272_),
    .C1(_09210_),
    .C2(_09465_),
    .ZN(_09686_));
 AND2_X1 _18988_ (.A1(_09684_),
    .A2(_09686_),
    .ZN(_09687_));
 AOI221_X1 _18989_ (.A(_09672_),
    .B1(_09677_),
    .B2(_09683_),
    .C1(_09687_),
    .C2(_09343_),
    .ZN(_09688_));
 AOI221_X1 _18990_ (.A(_09226_),
    .B1(_09206_),
    .B2(_09114_),
    .C1(_09332_),
    .C2(net123),
    .ZN(_09689_));
 OR3_X1 _18991_ (.A1(_09265_),
    .A2(_09377_),
    .A3(_09689_),
    .ZN(_09690_));
 OAI221_X1 _18992_ (.A(_09266_),
    .B1(_09325_),
    .B2(_09337_),
    .C1(_09113_),
    .C2(net122),
    .ZN(_09691_));
 NAND3_X1 _18993_ (.A1(_09489_),
    .A2(_09690_),
    .A3(_09691_),
    .ZN(_09692_));
 NOR4_X1 _18994_ (.A1(_09259_),
    .A2(_09449_),
    .A3(_09344_),
    .A4(_09345_),
    .ZN(_09693_));
 AND3_X1 _18995_ (.A1(_09241_),
    .A2(_09601_),
    .A3(_09305_),
    .ZN(_09694_));
 AOI211_X2 _18996_ (.A(_09058_),
    .B(_09328_),
    .C1(_09133_),
    .C2(net124),
    .ZN(_09695_));
 AOI21_X1 _18997_ (.A(_09063_),
    .B1(_09295_),
    .B2(_09269_),
    .ZN(_09696_));
 NOR3_X1 _18998_ (.A1(_09454_),
    .A2(_09695_),
    .A3(_09696_),
    .ZN(_09697_));
 NAND4_X1 _18999_ (.A1(_09203_),
    .A2(_09081_),
    .A3(_09123_),
    .A4(_09127_),
    .ZN(_09698_));
 OAI21_X1 _19000_ (.A(_09698_),
    .B1(_09247_),
    .B2(_14808_),
    .ZN(_09699_));
 MUX2_X1 _19001_ (.A(_09237_),
    .B(_09217_),
    .S(_09062_),
    .Z(_09700_));
 MUX2_X1 _19002_ (.A(_14822_),
    .B(_09700_),
    .S(_09133_),
    .Z(_09701_));
 OAI22_X2 _19003_ (.A1(_09387_),
    .A2(_09699_),
    .B1(_09701_),
    .B2(_09382_),
    .ZN(_09702_));
 OR4_X2 _19004_ (.A1(_09693_),
    .A2(_09702_),
    .A3(_09697_),
    .A4(_09694_),
    .ZN(_09703_));
 AOI22_X2 _19005_ (.A1(_09218_),
    .A2(_09216_),
    .B1(_09492_),
    .B2(_09256_),
    .ZN(_09704_));
 NAND4_X1 _19006_ (.A1(_09185_),
    .A2(_09309_),
    .A3(_09356_),
    .A4(_09704_),
    .ZN(_09705_));
 AOI21_X1 _19007_ (.A(_09521_),
    .B1(_09369_),
    .B2(_09646_),
    .ZN(_09706_));
 OAI21_X1 _19008_ (.A(_09705_),
    .B1(_09706_),
    .B2(_09185_),
    .ZN(_09707_));
 OAI221_X1 _19009_ (.A(_09692_),
    .B1(_09703_),
    .B2(_09080_),
    .C1(_09410_),
    .C2(_09707_),
    .ZN(_09708_));
 MUX2_X1 _19010_ (.A(_09688_),
    .B(_09708_),
    .S(_09246_),
    .Z(_00039_));
 INV_X1 _19011_ (.A(net1087),
    .ZN(_09709_));
 NOR2_X1 _19012_ (.A1(_09709_),
    .A2(_09102_),
    .ZN(_09710_));
 NOR2_X1 _19013_ (.A1(net1087),
    .A2(_09102_),
    .ZN(_09711_));
 BUF_X4 _19014_ (.A(\sa01_sr[7] ),
    .Z(_09712_));
 BUF_X16 clone127 (.A(_09727_),
    .Z(net610));
 XOR2_X2 _19016_ (.A(\sa11_sr[7] ),
    .B(_09712_),
    .Z(_09714_));
 BUF_X4 clone7 (.A(net124),
    .Z(net7));
 NOR2_X2 clone4 (.A1(net1227),
    .A2(_06449_),
    .ZN(net4));
 XNOR2_X2 _19019_ (.A(\sa21_sr[1] ),
    .B(\sa11_sr[1] ),
    .ZN(_09717_));
 XNOR2_X2 _19020_ (.A(net774),
    .B(_09714_),
    .ZN(_09718_));
 BUF_X4 _19021_ (.A(\sa01_sr[0] ),
    .Z(_09719_));
 BUF_X2 split138 (.A(_14970_),
    .Z(net138));
 NOR2_X4 clone174 (.A1(_13174_),
    .A2(net494),
    .ZN(net174));
 XOR2_X1 _19024_ (.A(\sa30_sub[1] ),
    .B(\sa11_sr[0] ),
    .Z(_09722_));
 XNOR2_X1 _19025_ (.A(_09722_),
    .B(_09719_),
    .ZN(_09723_));
 XNOR2_X2 _19026_ (.A(_09723_),
    .B(_09718_),
    .ZN(_09724_));
 MUX2_X2 _19027_ (.A(_09710_),
    .B(_09711_),
    .S(_09724_),
    .Z(_09725_));
 BUF_X32 _19028_ (.A(_08971_),
    .Z(_09726_));
 BUF_X32 _19029_ (.A(_09726_),
    .Z(_09727_));
 BUF_X32 _19030_ (.A(_09727_),
    .Z(_09728_));
 NAND3_X1 _19031_ (.A1(net1087),
    .A2(net610),
    .A3(_00443_),
    .ZN(_09729_));
 BUF_X8 _19032_ (.A(_09727_),
    .Z(_09730_));
 NAND2_X1 _19033_ (.A1(_09709_),
    .A2(_09730_),
    .ZN(_09731_));
 OAI21_X4 _19034_ (.A(_09729_),
    .B1(_09731_),
    .B2(_00443_),
    .ZN(_09732_));
 NOR2_X4 _19035_ (.A1(_09732_),
    .A2(_09725_),
    .ZN(_09733_));
 INV_X8 _19036_ (.A(_09733_),
    .ZN(_09734_));
 BUF_X16 _19037_ (.A(_09734_),
    .Z(_09735_));
 BUF_X32 _19038_ (.A(_09735_),
    .Z(_09736_));
 BUF_X32 _19039_ (.A(_09736_),
    .Z(_14832_));
 BUF_X4 clone12 (.A(_07426_),
    .Z(net12));
 BUF_X8 clone145 (.A(net720),
    .Z(net145));
 XNOR2_X2 _19042_ (.A(\sa11_sr[0] ),
    .B(net759),
    .ZN(_09739_));
 XNOR2_X1 _19043_ (.A(net642),
    .B(net669),
    .ZN(_09740_));
 NAND3_X1 _19044_ (.A1(net783),
    .A2(_09022_),
    .A3(_09714_),
    .ZN(_09741_));
 XNOR2_X2 _19045_ (.A(_09712_),
    .B(\sa11_sr[7] ),
    .ZN(_09742_));
 NOR2_X1 _19046_ (.A1(net782),
    .A2(_08992_),
    .ZN(_09743_));
 NAND2_X1 _19047_ (.A1(_09742_),
    .A2(_09743_),
    .ZN(_09744_));
 AOI21_X1 _19048_ (.A(_09740_),
    .B1(_09741_),
    .B2(_09744_),
    .ZN(_09745_));
 XOR2_X1 _19049_ (.A(net642),
    .B(net668),
    .Z(_09746_));
 NAND2_X1 _19050_ (.A1(_09714_),
    .A2(_09743_),
    .ZN(_09747_));
 NAND3_X1 _19051_ (.A1(net782),
    .A2(net948),
    .A3(_09742_),
    .ZN(_09748_));
 AOI21_X1 _19052_ (.A(_09746_),
    .B1(_09747_),
    .B2(_09748_),
    .ZN(_09749_));
 INV_X1 _19053_ (.A(net782),
    .ZN(_09750_));
 NAND3_X1 _19054_ (.A1(_09750_),
    .A2(_09726_),
    .A3(_00444_),
    .ZN(_09751_));
 NAND2_X1 _19055_ (.A1(net782),
    .A2(_09726_),
    .ZN(_09752_));
 OAI21_X1 _19056_ (.A(_09751_),
    .B1(_09752_),
    .B2(_00444_),
    .ZN(_09753_));
 OR3_X1 _19057_ (.A1(_09745_),
    .A2(_09749_),
    .A3(_09753_),
    .ZN(_09754_));
 BUF_X4 _19058_ (.A(_09754_),
    .Z(_09755_));
 INV_X16 _19059_ (.A(_09755_),
    .ZN(_09756_));
 BUF_X2 rebuffer134 (.A(_14829_),
    .Z(net617));
 BUF_X8 _19061_ (.A(_09756_),
    .Z(_14835_));
 INV_X2 clone173 (.A(net174),
    .ZN(net173));
 BUF_X4 _19063_ (.A(\sa30_sub[2] ),
    .Z(_09759_));
 XOR2_X2 _19064_ (.A(\sa11_sr[1] ),
    .B(_09759_),
    .Z(_09760_));
 XOR2_X1 _19065_ (.A(net752),
    .B(_09760_),
    .Z(_09761_));
 CLKBUF_X3 _19066_ (.A(\sa11_sr[2] ),
    .Z(_09762_));
 BUF_X4 _19067_ (.A(\sa21_sr[2] ),
    .Z(_09763_));
 XOR2_X2 _19068_ (.A(_09762_),
    .B(_09763_),
    .Z(_09764_));
 NAND3_X1 _19069_ (.A1(_06638_),
    .A2(net948),
    .A3(_09764_),
    .ZN(_09765_));
 XNOR2_X2 _19070_ (.A(_09762_),
    .B(_09763_),
    .ZN(_09766_));
 NOR2_X1 _19071_ (.A1(_06638_),
    .A2(_08971_),
    .ZN(_09767_));
 NAND2_X1 _19072_ (.A1(_09766_),
    .A2(_09767_),
    .ZN(_09768_));
 AOI21_X2 _19073_ (.A(_09761_),
    .B1(_09765_),
    .B2(_09768_),
    .ZN(_09769_));
 XNOR2_X1 _19074_ (.A(net752),
    .B(_09760_),
    .ZN(_09770_));
 NAND2_X1 _19075_ (.A1(_09764_),
    .A2(_09767_),
    .ZN(_09771_));
 NAND3_X1 _19076_ (.A1(_06638_),
    .A2(_09010_),
    .A3(_09766_),
    .ZN(_09772_));
 AOI21_X2 _19077_ (.A(_09770_),
    .B1(_09771_),
    .B2(_09772_),
    .ZN(_09773_));
 INV_X1 _19078_ (.A(_06638_),
    .ZN(_09774_));
 NAND3_X1 _19079_ (.A1(_09774_),
    .A2(_08972_),
    .A3(_00445_),
    .ZN(_09775_));
 NAND2_X1 _19080_ (.A1(_06638_),
    .A2(_08972_),
    .ZN(_09776_));
 OAI21_X2 _19081_ (.A(_09775_),
    .B1(_09776_),
    .B2(_00445_),
    .ZN(_09777_));
 NOR3_X4 _19082_ (.A1(_09769_),
    .A2(_09773_),
    .A3(_09777_),
    .ZN(_09778_));
 INV_X8 _19083_ (.A(_09778_),
    .ZN(_09779_));
 BUF_X4 _19084_ (.A(_09779_),
    .Z(_09780_));
 BUF_X4 _19085_ (.A(_09780_),
    .Z(_09781_));
 BUF_X4 _19086_ (.A(_09781_),
    .Z(_09782_));
 BUF_X4 _19087_ (.A(_09782_),
    .Z(_14851_));
 BUF_X4 _19088_ (.A(_09755_),
    .Z(_14826_));
 BUF_X4 _19089_ (.A(_09778_),
    .Z(_09783_));
 BUF_X4 _19090_ (.A(_09783_),
    .Z(_09784_));
 BUF_X4 _19091_ (.A(_09784_),
    .Z(_14844_));
 BUF_X2 _19092_ (.A(\sa11_sr[5] ),
    .Z(_09785_));
 CLKBUF_X3 _19093_ (.A(\sa11_sr[6] ),
    .Z(_09786_));
 BUF_X4 _19094_ (.A(\sa21_sr[6] ),
    .Z(_09787_));
 XNOR2_X2 _19095_ (.A(_09786_),
    .B(_09787_),
    .ZN(_09788_));
 CLKBUF_X3 _19096_ (.A(\sa01_sr[5] ),
    .Z(_09789_));
 CLKBUF_X3 _19097_ (.A(\sa30_sub[6] ),
    .Z(_09790_));
 XNOR2_X1 _19098_ (.A(_09789_),
    .B(_09790_),
    .ZN(_09791_));
 XNOR2_X1 _19099_ (.A(_09788_),
    .B(_09791_),
    .ZN(_09792_));
 XNOR2_X1 _19100_ (.A(_09785_),
    .B(_09792_),
    .ZN(_09793_));
 MUX2_X2 _19101_ (.A(\text_in_r[94] ),
    .B(_09793_),
    .S(_09074_),
    .Z(_09794_));
 XOR2_X2 _19102_ (.A(_06697_),
    .B(_09794_),
    .Z(_09795_));
 BUF_X4 _19103_ (.A(\sa21_sr[7] ),
    .Z(_09796_));
 XNOR2_X2 _19104_ (.A(net705),
    .B(_09796_),
    .ZN(_09797_));
 BUF_X2 _19105_ (.A(\sa01_sr[6] ),
    .Z(_09798_));
 BUF_X8 _19106_ (.A(\sa30_sub[7] ),
    .Z(_09799_));
 XNOR2_X1 _19107_ (.A(_09798_),
    .B(_09799_),
    .ZN(_09800_));
 XNOR2_X1 _19108_ (.A(net667),
    .B(_09800_),
    .ZN(_09801_));
 XNOR2_X1 _19109_ (.A(_09786_),
    .B(_09801_),
    .ZN(_09802_));
 BUF_X4 _19110_ (.A(_09138_),
    .Z(_09803_));
 MUX2_X1 _19111_ (.A(\text_in_r[95] ),
    .B(_09802_),
    .S(_09803_),
    .Z(_09804_));
 XNOR2_X2 _19112_ (.A(_06711_),
    .B(_09804_),
    .ZN(_09805_));
 NOR2_X4 _19113_ (.A1(_09795_),
    .A2(_09805_),
    .ZN(_09806_));
 INV_X1 _19114_ (.A(_06688_),
    .ZN(_09807_));
 CLKBUF_X3 _19115_ (.A(\sa11_sr[4] ),
    .Z(_09808_));
 CLKBUF_X3 _19116_ (.A(\sa30_sub[5] ),
    .Z(_09809_));
 XNOR2_X1 _19117_ (.A(_09808_),
    .B(_09809_),
    .ZN(_09810_));
 NOR3_X1 _19118_ (.A1(_09807_),
    .A2(_09180_),
    .A3(_09810_),
    .ZN(_09811_));
 NOR3_X1 _19119_ (.A1(_06688_),
    .A2(_09180_),
    .A3(_09810_),
    .ZN(_09812_));
 BUF_X2 _19120_ (.A(\sa01_sr[4] ),
    .Z(_09813_));
 BUF_X4 _19121_ (.A(\sa21_sr[5] ),
    .Z(_09814_));
 XNOR2_X1 _19122_ (.A(_09785_),
    .B(_09814_),
    .ZN(_09815_));
 XNOR2_X2 _19123_ (.A(_09813_),
    .B(_09815_),
    .ZN(_09816_));
 MUX2_X1 _19124_ (.A(_09811_),
    .B(_09812_),
    .S(_09816_),
    .Z(_09817_));
 BUF_X32 _19125_ (.A(_09728_),
    .Z(_09818_));
 XOR2_X2 _19126_ (.A(_09808_),
    .B(_09809_),
    .Z(_09819_));
 NOR3_X1 _19127_ (.A1(_06688_),
    .A2(net582),
    .A3(_09819_),
    .ZN(_09820_));
 NOR3_X1 _19128_ (.A1(_09807_),
    .A2(net582),
    .A3(_09819_),
    .ZN(_09821_));
 MUX2_X1 _19129_ (.A(_09820_),
    .B(_09821_),
    .S(_09816_),
    .Z(_09822_));
 BUF_X16 _19130_ (.A(_08974_),
    .Z(_09823_));
 BUF_X8 _19131_ (.A(_09823_),
    .Z(_09824_));
 NAND3_X1 _19132_ (.A1(_06688_),
    .A2(_09824_),
    .A3(\text_in_r[93] ),
    .ZN(_09825_));
 NAND2_X1 _19133_ (.A1(_09807_),
    .A2(_09824_),
    .ZN(_09826_));
 OAI21_X2 _19134_ (.A(_09825_),
    .B1(_09826_),
    .B2(\text_in_r[93] ),
    .ZN(_09827_));
 NOR3_X4 _19135_ (.A1(_09817_),
    .A2(_09822_),
    .A3(_09827_),
    .ZN(_09828_));
 BUF_X4 _19136_ (.A(_09828_),
    .Z(_09829_));
 CLKBUF_X3 _19137_ (.A(_09829_),
    .Z(_09830_));
 BUF_X4 _19138_ (.A(_09779_),
    .Z(_09831_));
 NOR2_X1 _19139_ (.A1(_06657_),
    .A2(_08973_),
    .ZN(_09832_));
 INV_X1 _19140_ (.A(_06657_),
    .ZN(_09833_));
 NOR2_X1 _19141_ (.A1(_09833_),
    .A2(_08973_),
    .ZN(_09834_));
 BUF_X4 _19142_ (.A(\sa01_sr[2] ),
    .Z(_09835_));
 BUF_X4 _19143_ (.A(\sa21_sr[3] ),
    .Z(_09836_));
 XNOR2_X1 _19144_ (.A(_09835_),
    .B(_09836_),
    .ZN(_09837_));
 XNOR2_X2 _19145_ (.A(_09712_),
    .B(_09837_),
    .ZN(_09838_));
 CLKBUF_X3 _19146_ (.A(\sa11_sr[3] ),
    .Z(_09839_));
 XOR2_X2 _19147_ (.A(\sa11_sr[7] ),
    .B(_09839_),
    .Z(_09840_));
 CLKBUF_X3 _19148_ (.A(\sa30_sub[3] ),
    .Z(_09841_));
 XNOR2_X1 _19149_ (.A(_09762_),
    .B(_09841_),
    .ZN(_09842_));
 XNOR2_X1 _19150_ (.A(_09840_),
    .B(_09842_),
    .ZN(_09843_));
 XNOR2_X1 _19151_ (.A(_09838_),
    .B(_09843_),
    .ZN(_09844_));
 MUX2_X1 _19152_ (.A(_09832_),
    .B(_09834_),
    .S(_09844_),
    .Z(_09845_));
 BUF_X4 _19153_ (.A(_09845_),
    .Z(_09846_));
 OR3_X2 _19154_ (.A1(_09833_),
    .A2(_09074_),
    .A3(\text_in_r[91] ),
    .ZN(_09847_));
 NAND3_X2 _19155_ (.A1(_09833_),
    .A2(_08994_),
    .A3(\text_in_r[91] ),
    .ZN(_09848_));
 NAND2_X4 _19156_ (.A1(_09847_),
    .A2(_09848_),
    .ZN(_09849_));
 NOR2_X1 _19157_ (.A1(_09846_),
    .A2(_09849_),
    .ZN(_09850_));
 BUF_X4 _19158_ (.A(_09850_),
    .Z(_09851_));
 BUF_X8 _19159_ (.A(_09851_),
    .Z(_09852_));
 BUF_X8 _19160_ (.A(_14830_),
    .Z(_09853_));
 INV_X4 _19161_ (.A(_09853_),
    .ZN(_09854_));
 NAND2_X1 _19162_ (.A1(_09833_),
    .A2(net594),
    .ZN(_09855_));
 BUF_X32 _19163_ (.A(_09099_),
    .Z(_09856_));
 NAND2_X1 _19164_ (.A1(_06657_),
    .A2(net1085),
    .ZN(_09857_));
 MUX2_X2 _19165_ (.A(_09855_),
    .B(_09857_),
    .S(_09844_),
    .Z(_09858_));
 BUF_X8 _19166_ (.A(_09858_),
    .Z(_09859_));
 AND2_X2 _19167_ (.A1(_09847_),
    .A2(_09848_),
    .ZN(_09860_));
 BUF_X8 _19168_ (.A(_09860_),
    .Z(_09861_));
 AOI21_X4 _19169_ (.A(_09756_),
    .B1(_09859_),
    .B2(_09861_),
    .ZN(_09862_));
 BUF_X4 _19170_ (.A(_09735_),
    .Z(_09863_));
 AOI221_X2 _19171_ (.A(_09831_),
    .B1(_09852_),
    .B2(_09854_),
    .C1(_09862_),
    .C2(_09863_),
    .ZN(_09864_));
 INV_X1 _19172_ (.A(_06673_),
    .ZN(_09865_));
 NOR2_X1 _19173_ (.A1(_09865_),
    .A2(_09818_),
    .ZN(_09866_));
 NOR2_X1 _19174_ (.A1(_06673_),
    .A2(_09818_),
    .ZN(_09867_));
 CLKBUF_X3 _19175_ (.A(\sa01_sr[3] ),
    .Z(_09868_));
 BUF_X4 _19176_ (.A(\sa21_sr[4] ),
    .Z(_09869_));
 XNOR2_X1 _19177_ (.A(_09868_),
    .B(_09869_),
    .ZN(_09870_));
 XNOR2_X1 _19178_ (.A(_09712_),
    .B(_09870_),
    .ZN(_09871_));
 BUF_X4 _19179_ (.A(\sa30_sub[4] ),
    .Z(_09872_));
 XOR2_X1 _19180_ (.A(_09808_),
    .B(_09872_),
    .Z(_09873_));
 XNOR2_X1 _19181_ (.A(_09840_),
    .B(_09873_),
    .ZN(_09874_));
 XNOR2_X1 _19182_ (.A(_09871_),
    .B(_09874_),
    .ZN(_09875_));
 MUX2_X2 _19183_ (.A(_09866_),
    .B(_09867_),
    .S(_09875_),
    .Z(_09876_));
 NAND3_X1 _19184_ (.A1(_09865_),
    .A2(_08996_),
    .A3(\text_in_r[92] ),
    .ZN(_09877_));
 NAND2_X1 _19185_ (.A1(_06673_),
    .A2(_09135_),
    .ZN(_09878_));
 OAI21_X4 _19186_ (.A(_09877_),
    .B1(_09878_),
    .B2(\text_in_r[92] ),
    .ZN(_09879_));
 NOR2_X4 _19187_ (.A1(_09876_),
    .A2(_09879_),
    .ZN(_09880_));
 BUF_X4 _19188_ (.A(_09880_),
    .Z(_09881_));
 OAI21_X4 _19189_ (.A(_09779_),
    .B1(_09846_),
    .B2(_09849_),
    .ZN(_09882_));
 BUF_X1 split160 (.A(_15268_),
    .Z(net160));
 INV_X2 _19191_ (.A(net619),
    .ZN(_09884_));
 OAI21_X1 _19192_ (.A(_09881_),
    .B1(_09882_),
    .B2(_09884_),
    .ZN(_09885_));
 NAND2_X4 _19193_ (.A1(_09859_),
    .A2(_09861_),
    .ZN(_09886_));
 NOR3_X4 _19194_ (.A1(_09756_),
    .A2(_09846_),
    .A3(_09849_),
    .ZN(_09887_));
 AOI221_X2 _19195_ (.A(_09780_),
    .B1(_09886_),
    .B2(_09854_),
    .C1(_09887_),
    .C2(_09735_),
    .ZN(_09888_));
 OR2_X2 _19196_ (.A1(_09876_),
    .A2(_09879_),
    .ZN(_09889_));
 BUF_X4 _19197_ (.A(_09889_),
    .Z(_09890_));
 BUF_X4 _19198_ (.A(_09890_),
    .Z(_09891_));
 NAND3_X2 _19199_ (.A1(_09779_),
    .A2(_09859_),
    .A3(_09861_),
    .ZN(_09892_));
 CLKBUF_X3 _19200_ (.A(_09892_),
    .Z(_09893_));
 BUF_X4 _19201_ (.A(_14836_),
    .Z(_09894_));
 OAI21_X1 _19202_ (.A(_09891_),
    .B1(_09893_),
    .B2(_09894_),
    .ZN(_09895_));
 OAI221_X1 _19203_ (.A(_09830_),
    .B1(_09864_),
    .B2(_09885_),
    .C1(_09888_),
    .C2(_09895_),
    .ZN(_09896_));
 BUF_X4 _19204_ (.A(_09886_),
    .Z(_09897_));
 NOR3_X4 _19205_ (.A1(_09778_),
    .A2(_09846_),
    .A3(_09849_),
    .ZN(_09898_));
 BUF_X4 clone15 (.A(_07377_),
    .Z(net15));
 BUF_X4 _19207_ (.A(net485),
    .Z(_09900_));
 AOI221_X1 _19208_ (.A(_09880_),
    .B1(_09897_),
    .B2(_14849_),
    .C1(_09898_),
    .C2(_09900_),
    .ZN(_09901_));
 OR2_X1 _19209_ (.A1(_09830_),
    .A2(_09901_),
    .ZN(_09902_));
 BUF_X4 _19210_ (.A(_09890_),
    .Z(_09903_));
 BUF_X4 _19211_ (.A(_09903_),
    .Z(_09904_));
 NOR2_X4 _19212_ (.A1(_09756_),
    .A2(_09779_),
    .ZN(_09905_));
 BUF_X2 clone144 (.A(_02278_),
    .Z(net144));
 INV_X4 _19214_ (.A(_14833_),
    .ZN(_09907_));
 AOI221_X2 _19215_ (.A(_09886_),
    .B1(_09905_),
    .B2(_09734_),
    .C1(_09907_),
    .C2(_09779_),
    .ZN(_09908_));
 BUF_X4 _19216_ (.A(_14828_),
    .Z(_09909_));
 BUF_X4 _19217_ (.A(_09846_),
    .Z(_09910_));
 BUF_X4 _19218_ (.A(_09849_),
    .Z(_09911_));
 OAI21_X2 _19219_ (.A(_09783_),
    .B1(_09910_),
    .B2(_09911_),
    .ZN(_09912_));
 NOR2_X1 _19220_ (.A1(_09909_),
    .A2(_09912_),
    .ZN(_09913_));
 BUF_X4 _19221_ (.A(_09859_),
    .Z(_09914_));
 BUF_X4 _19222_ (.A(_09861_),
    .Z(_09915_));
 NAND3_X2 _19223_ (.A1(_09853_),
    .A2(_09914_),
    .A3(_09915_),
    .ZN(_09916_));
 OAI21_X4 _19224_ (.A(_09756_),
    .B1(_09910_),
    .B2(_09911_),
    .ZN(_09917_));
 AOI21_X1 _19225_ (.A(_09784_),
    .B1(_09916_),
    .B2(_09917_),
    .ZN(_09918_));
 NOR4_X2 _19226_ (.A1(_09904_),
    .A2(_09908_),
    .A3(_09913_),
    .A4(_09918_),
    .ZN(_09919_));
 OAI21_X1 _19227_ (.A(_09896_),
    .B1(_09919_),
    .B2(_09902_),
    .ZN(_09920_));
 AND2_X2 _19228_ (.A1(_09806_),
    .A2(_09920_),
    .ZN(_09921_));
 BUF_X4 _19229_ (.A(_09881_),
    .Z(_09922_));
 BUF_X4 _19230_ (.A(_09795_),
    .Z(_09923_));
 CLKBUF_X3 _19231_ (.A(_09852_),
    .Z(_09924_));
 NOR2_X1 _19232_ (.A1(net113),
    .A2(_09924_),
    .ZN(_09925_));
 NAND2_X1 _19233_ (.A1(_09755_),
    .A2(_09780_),
    .ZN(_09926_));
 CLKBUF_X3 _19234_ (.A(_09912_),
    .Z(_09927_));
 BUF_X8 _19235_ (.A(net707),
    .Z(_09928_));
 OAI221_X1 _19236_ (.A(_09923_),
    .B1(_09925_),
    .B2(_09926_),
    .C1(_09927_),
    .C2(_09928_),
    .ZN(_09929_));
 XNOR2_X2 _19237_ (.A(_06697_),
    .B(_09794_),
    .ZN(_09930_));
 BUF_X4 _19238_ (.A(_09930_),
    .Z(_09931_));
 CLKBUF_X3 _19239_ (.A(_09851_),
    .Z(_09932_));
 OAI21_X4 _19240_ (.A(_09756_),
    .B1(_09732_),
    .B2(_09725_),
    .ZN(_09933_));
 AND2_X1 _19241_ (.A1(_09932_),
    .A2(_09933_),
    .ZN(_09934_));
 CLKBUF_X3 _19242_ (.A(_09831_),
    .Z(_09935_));
 OAI21_X1 _19243_ (.A(_09935_),
    .B1(_09924_),
    .B2(_09909_),
    .ZN(_09936_));
 NAND3_X4 _19244_ (.A1(net486),
    .A2(_09859_),
    .A3(_09861_),
    .ZN(_09937_));
 BUF_X4 _19245_ (.A(_09852_),
    .Z(_09938_));
 OAI21_X1 _19246_ (.A(_09937_),
    .B1(_09938_),
    .B2(_09894_),
    .ZN(_09939_));
 CLKBUF_X3 _19247_ (.A(_09781_),
    .Z(_09940_));
 OAI221_X1 _19248_ (.A(_09931_),
    .B1(_09934_),
    .B2(_09936_),
    .C1(_09939_),
    .C2(_09940_),
    .ZN(_09941_));
 AND3_X1 _19249_ (.A1(_09922_),
    .A2(_09929_),
    .A3(_09941_),
    .ZN(_09942_));
 BUF_X4 _19250_ (.A(_09863_),
    .Z(_09943_));
 OAI21_X4 _19251_ (.A(_09755_),
    .B1(_09910_),
    .B2(_09911_),
    .ZN(_09944_));
 MUX2_X1 _19252_ (.A(_09893_),
    .B(_09944_),
    .S(_09930_),
    .Z(_09945_));
 NOR2_X1 _19253_ (.A1(_09943_),
    .A2(_09945_),
    .ZN(_09946_));
 NAND3_X4 _19254_ (.A1(_09756_),
    .A2(_09914_),
    .A3(_09915_),
    .ZN(_09947_));
 BUF_X4 _19255_ (.A(_09783_),
    .Z(_09948_));
 BUF_X4 _19256_ (.A(_09948_),
    .Z(_09949_));
 AOI21_X1 _19257_ (.A(_09947_),
    .B1(_09931_),
    .B2(_09949_),
    .ZN(_09950_));
 BUF_X4 _19258_ (.A(_09897_),
    .Z(_09951_));
 BUF_X4 clone107 (.A(net935),
    .Z(net107));
 MUX2_X1 _19260_ (.A(net111),
    .B(_14842_),
    .S(_09780_),
    .Z(_09953_));
 NAND3_X1 _19261_ (.A1(_09795_),
    .A2(_09953_),
    .A3(_09951_),
    .ZN(_09954_));
 NOR2_X4 _19262_ (.A1(_09755_),
    .A2(_09780_),
    .ZN(_09955_));
 AOI22_X1 _19263_ (.A1(_09863_),
    .A2(_09887_),
    .B1(_09955_),
    .B2(_09951_),
    .ZN(_09956_));
 OAI21_X1 _19264_ (.A(_09954_),
    .B1(_09956_),
    .B2(_09795_),
    .ZN(_09957_));
 NOR4_X2 _19265_ (.A1(_09957_),
    .A2(_09922_),
    .A3(_09950_),
    .A4(_09946_),
    .ZN(_09958_));
 CLKBUF_X3 _19266_ (.A(_09805_),
    .Z(_09959_));
 NAND2_X1 _19267_ (.A1(_09959_),
    .A2(_09830_),
    .ZN(_09960_));
 NOR3_X1 _19268_ (.A1(_09958_),
    .A2(_09942_),
    .A3(_09960_),
    .ZN(_09961_));
 NOR2_X1 _19269_ (.A1(_09930_),
    .A2(_09805_),
    .ZN(_09962_));
 BUF_X4 _19270_ (.A(_09880_),
    .Z(_09963_));
 NAND2_X1 _19271_ (.A1(_09780_),
    .A2(net485),
    .ZN(_09964_));
 OAI21_X4 _19272_ (.A(_09778_),
    .B1(_09732_),
    .B2(net567),
    .ZN(_09965_));
 NAND3_X1 _19273_ (.A1(_09852_),
    .A2(_09964_),
    .A3(_09965_),
    .ZN(_09966_));
 NAND2_X1 _19274_ (.A1(_09963_),
    .A2(_09966_),
    .ZN(_09967_));
 INV_X2 _19275_ (.A(_09894_),
    .ZN(_09968_));
 AOI21_X1 _19276_ (.A(_09955_),
    .B1(_09831_),
    .B2(_09968_),
    .ZN(_09969_));
 OAI21_X1 _19277_ (.A(_09828_),
    .B1(_09932_),
    .B2(_09969_),
    .ZN(_09970_));
 OAI21_X1 _19278_ (.A(_09962_),
    .B1(_09967_),
    .B2(_09970_),
    .ZN(_09971_));
 NOR2_X1 _19279_ (.A1(_09755_),
    .A2(_09882_),
    .ZN(_09972_));
 AOI21_X4 _19280_ (.A(_09779_),
    .B1(_09858_),
    .B2(_09860_),
    .ZN(_09973_));
 AOI221_X2 _19281_ (.A(_09972_),
    .B1(_09933_),
    .B2(_09973_),
    .C1(_09928_),
    .C2(_09898_),
    .ZN(_09974_));
 NOR2_X1 _19282_ (.A1(_09829_),
    .A2(_09903_),
    .ZN(_09975_));
 INV_X2 _19283_ (.A(_09909_),
    .ZN(_09976_));
 NAND3_X4 _19284_ (.A1(_09778_),
    .A2(_09859_),
    .A3(_09861_),
    .ZN(_09977_));
 OAI222_X2 _19285_ (.A1(_09928_),
    .A2(_09912_),
    .B1(_09892_),
    .B2(_09976_),
    .C1(_09977_),
    .C2(_09853_),
    .ZN(_09978_));
 OAI21_X4 _19286_ (.A(net111),
    .B1(_09910_),
    .B2(_09911_),
    .ZN(_09979_));
 NAND3_X2 _19287_ (.A1(net618),
    .A2(_09914_),
    .A3(_09915_),
    .ZN(_09980_));
 NAND3_X1 _19288_ (.A1(_09783_),
    .A2(_09979_),
    .A3(_09980_),
    .ZN(_09981_));
 OAI21_X1 _19289_ (.A(_09981_),
    .B1(_09893_),
    .B2(_09928_),
    .ZN(_09982_));
 OR3_X2 _19290_ (.A1(_09817_),
    .A2(_09822_),
    .A3(_09827_),
    .ZN(_09983_));
 BUF_X4 _19291_ (.A(_09983_),
    .Z(_09984_));
 MUX2_X1 _19292_ (.A(_09978_),
    .B(_09982_),
    .S(_09984_),
    .Z(_09985_));
 AOI221_X1 _19293_ (.A(_09971_),
    .B1(_09974_),
    .B2(_09975_),
    .C1(_09985_),
    .C2(_09904_),
    .ZN(_09986_));
 NAND2_X1 _19294_ (.A1(_09882_),
    .A2(_09977_),
    .ZN(_09987_));
 NAND2_X1 _19295_ (.A1(_09909_),
    .A2(_09987_),
    .ZN(_09988_));
 INV_X4 _19296_ (.A(net617),
    .ZN(_09989_));
 AOI221_X2 _19297_ (.A(_09795_),
    .B1(_09973_),
    .B2(_09989_),
    .C1(_09898_),
    .C2(_14836_),
    .ZN(_09990_));
 NOR3_X4 _19298_ (.A1(_09779_),
    .A2(_09846_),
    .A3(_09849_),
    .ZN(_09991_));
 NAND2_X4 _19299_ (.A1(_09756_),
    .A2(_09778_),
    .ZN(_09992_));
 OAI21_X1 _19300_ (.A(_09892_),
    .B1(_09992_),
    .B2(_09850_),
    .ZN(_09993_));
 AOI222_X2 _19301_ (.A1(_09854_),
    .A2(_09991_),
    .B1(_09993_),
    .B2(_09734_),
    .C1(_09779_),
    .C2(_09862_),
    .ZN(_09994_));
 AOI221_X2 _19302_ (.A(_09890_),
    .B1(_09988_),
    .B2(_09990_),
    .C1(_09994_),
    .C2(_09795_),
    .ZN(_09995_));
 BUF_X4 _19303_ (.A(_09984_),
    .Z(_09996_));
 NAND2_X1 _19304_ (.A1(_09805_),
    .A2(_09996_),
    .ZN(_09997_));
 MUX2_X1 _19305_ (.A(_14842_),
    .B(_09735_),
    .S(_09851_),
    .Z(_09998_));
 NOR2_X2 _19306_ (.A1(net112),
    .A2(_09897_),
    .ZN(_09999_));
 OAI22_X1 _19307_ (.A1(_09781_),
    .A2(_09998_),
    .B1(_09999_),
    .B2(_09926_),
    .ZN(_10000_));
 AOI21_X1 _19308_ (.A(_09937_),
    .B1(_09831_),
    .B2(_09733_),
    .ZN(_10001_));
 NOR2_X1 _19309_ (.A1(_09900_),
    .A2(_09783_),
    .ZN(_10002_));
 BUF_X8 _19310_ (.A(net936),
    .Z(_10003_));
 NAND2_X1 _19311_ (.A1(net934),
    .A2(_09852_),
    .ZN(_10004_));
 AOI21_X1 _19312_ (.A(_10001_),
    .B1(_10002_),
    .B2(_10004_),
    .ZN(_10005_));
 MUX2_X1 _19313_ (.A(_10000_),
    .B(_10005_),
    .S(_09930_),
    .Z(_10006_));
 AOI211_X2 _19314_ (.A(_09995_),
    .B(_09997_),
    .C1(_10006_),
    .C2(_09904_),
    .ZN(_10007_));
 OR4_X4 _19315_ (.A1(_09961_),
    .A2(_10007_),
    .A3(_09986_),
    .A4(_09921_),
    .ZN(_00040_));
 NOR2_X2 _19316_ (.A1(_09984_),
    .A2(_09963_),
    .ZN(_10008_));
 BUF_X4 rebuffer370 (.A(_11130_),
    .Z(net883));
 OAI21_X1 _19318_ (.A(_10008_),
    .B1(_09947_),
    .B2(net108),
    .ZN(_10009_));
 INV_X2 _19319_ (.A(_14842_),
    .ZN(_10010_));
 NOR2_X1 _19320_ (.A1(_10010_),
    .A2(_09932_),
    .ZN(_10011_));
 OAI22_X1 _19321_ (.A1(net113),
    .A2(_09927_),
    .B1(_10011_),
    .B2(_09949_),
    .ZN(_10012_));
 OAI21_X4 _19322_ (.A(_09989_),
    .B1(_09910_),
    .B2(_09911_),
    .ZN(_10013_));
 NAND3_X2 _19323_ (.A1(_09976_),
    .A2(_09914_),
    .A3(_09915_),
    .ZN(_10014_));
 AOI21_X1 _19324_ (.A(_09935_),
    .B1(_10013_),
    .B2(_10014_),
    .ZN(_10015_));
 OAI21_X4 _19325_ (.A(net707),
    .B1(_09910_),
    .B2(_09911_),
    .ZN(_10016_));
 AOI21_X1 _19326_ (.A(_09949_),
    .B1(_09947_),
    .B2(_10016_),
    .ZN(_10017_));
 NOR2_X1 _19327_ (.A1(_10015_),
    .A2(_10017_),
    .ZN(_10018_));
 NAND2_X1 _19328_ (.A1(_09996_),
    .A2(_09891_),
    .ZN(_10019_));
 OAI221_X1 _19329_ (.A(_09962_),
    .B1(_10009_),
    .B2(_10012_),
    .C1(_10018_),
    .C2(_10019_),
    .ZN(_10020_));
 NOR2_X1 _19330_ (.A1(_09907_),
    .A2(_09951_),
    .ZN(_10021_));
 NAND2_X4 _19331_ (.A1(_10013_),
    .A2(_09784_),
    .ZN(_10022_));
 BUF_X4 _19332_ (.A(_09897_),
    .Z(_10023_));
 AND2_X1 _19333_ (.A1(_10023_),
    .A2(_09933_),
    .ZN(_10024_));
 BUF_X4 _19334_ (.A(_09784_),
    .Z(_10025_));
 OAI221_X1 _19335_ (.A(_09830_),
    .B1(_10021_),
    .B2(_10022_),
    .C1(_10024_),
    .C2(_10025_),
    .ZN(_10026_));
 AOI21_X4 _19336_ (.A(_09755_),
    .B1(_09859_),
    .B2(_09861_),
    .ZN(_10027_));
 AOI22_X1 _19337_ (.A1(net108),
    .A2(_10027_),
    .B1(_09898_),
    .B2(net110),
    .ZN(_10028_));
 AOI21_X4 _19338_ (.A(_09783_),
    .B1(_09914_),
    .B2(_09915_),
    .ZN(_10029_));
 NOR2_X2 _19339_ (.A1(_10029_),
    .A2(_09991_),
    .ZN(_10030_));
 OAI21_X1 _19340_ (.A(_10028_),
    .B1(_10030_),
    .B2(_14835_),
    .ZN(_10031_));
 BUF_X4 _19341_ (.A(_09828_),
    .Z(_10032_));
 CLKBUF_X3 _19342_ (.A(_10032_),
    .Z(_10033_));
 OAI21_X1 _19343_ (.A(_10026_),
    .B1(_10031_),
    .B2(_10033_),
    .ZN(_10034_));
 BUF_X4 _19344_ (.A(_09881_),
    .Z(_10035_));
 AOI21_X1 _19345_ (.A(_10020_),
    .B1(_10034_),
    .B2(_10035_),
    .ZN(_10036_));
 INV_X2 _19346_ (.A(_09805_),
    .ZN(_10037_));
 NAND3_X2 _19347_ (.A1(_09854_),
    .A2(_09914_),
    .A3(_09915_),
    .ZN(_10038_));
 NAND2_X1 _19348_ (.A1(net112),
    .A2(_10027_),
    .ZN(_10039_));
 AOI21_X1 _19349_ (.A(_10025_),
    .B1(_10038_),
    .B2(_10039_),
    .ZN(_10040_));
 AOI21_X2 _19350_ (.A(_09900_),
    .B1(_09914_),
    .B2(_09915_),
    .ZN(_10041_));
 NOR2_X1 _19351_ (.A1(_09935_),
    .A2(_10041_),
    .ZN(_10042_));
 NAND3_X4 _19352_ (.A1(net536),
    .A2(_09859_),
    .A3(_09861_),
    .ZN(_10043_));
 AND2_X1 _19353_ (.A1(_10042_),
    .A2(net645),
    .ZN(_10044_));
 OAI21_X1 _19354_ (.A(_09996_),
    .B1(_10040_),
    .B2(_10044_),
    .ZN(_10045_));
 NAND2_X1 _19355_ (.A1(_09923_),
    .A2(_09891_),
    .ZN(_10046_));
 NAND3_X1 _19356_ (.A1(_09782_),
    .A2(_09947_),
    .A3(_09979_),
    .ZN(_10047_));
 OAI21_X1 _19357_ (.A(_09916_),
    .B1(_09938_),
    .B2(net878),
    .ZN(_10048_));
 CLKBUF_X3 _19358_ (.A(_09935_),
    .Z(_10049_));
 OAI21_X1 _19359_ (.A(_10047_),
    .B1(_10048_),
    .B2(_10049_),
    .ZN(_10050_));
 AOI21_X1 _19360_ (.A(_10046_),
    .B1(_10050_),
    .B2(_09830_),
    .ZN(_10051_));
 AOI21_X1 _19361_ (.A(_10037_),
    .B1(_10045_),
    .B2(_10051_),
    .ZN(_10052_));
 AOI21_X2 _19362_ (.A(_09907_),
    .B1(_09859_),
    .B2(_09861_),
    .ZN(_10053_));
 NOR3_X2 _19363_ (.A1(_10053_),
    .A2(_09887_),
    .A3(_09780_),
    .ZN(_10054_));
 XNOR2_X1 _19364_ (.A(_09735_),
    .B(_09851_),
    .ZN(_10055_));
 AOI211_X2 _19365_ (.A(_09828_),
    .B(_10054_),
    .C1(_10055_),
    .C2(_09781_),
    .ZN(_10056_));
 XNOR2_X2 _19366_ (.A(_09756_),
    .B(_09780_),
    .ZN(_10057_));
 NOR3_X1 _19367_ (.A1(net107),
    .A2(_09932_),
    .A3(_10057_),
    .ZN(_10058_));
 MUX2_X1 _19368_ (.A(_09976_),
    .B(_09756_),
    .S(_09783_),
    .Z(_10059_));
 OAI21_X1 _19369_ (.A(_09828_),
    .B1(_09951_),
    .B2(_10059_),
    .ZN(_10060_));
 OAI21_X1 _19370_ (.A(_09903_),
    .B1(_10058_),
    .B2(_10060_),
    .ZN(_10061_));
 NOR2_X1 _19371_ (.A1(_09935_),
    .A2(_09933_),
    .ZN(_10062_));
 OAI21_X1 _19372_ (.A(_09932_),
    .B1(_09784_),
    .B2(_09968_),
    .ZN(_10063_));
 OAI21_X1 _19373_ (.A(_09881_),
    .B1(_10062_),
    .B2(_10063_),
    .ZN(_10064_));
 NOR3_X1 _19374_ (.A1(_14852_),
    .A2(_10032_),
    .A3(_09938_),
    .ZN(_10065_));
 OAI221_X1 _19375_ (.A(_09931_),
    .B1(_10061_),
    .B2(_10056_),
    .C1(_10064_),
    .C2(_10065_),
    .ZN(_10066_));
 NOR2_X1 _19376_ (.A1(_09930_),
    .A2(_09903_),
    .ZN(_10067_));
 MUX2_X1 _19377_ (.A(_09907_),
    .B(_09733_),
    .S(_09780_),
    .Z(_10068_));
 OAI21_X1 _19378_ (.A(_10032_),
    .B1(_09938_),
    .B2(_10068_),
    .ZN(_10069_));
 NAND2_X1 _19379_ (.A1(_09909_),
    .A2(_09779_),
    .ZN(_10070_));
 NOR2_X1 _19380_ (.A1(_09897_),
    .A2(_09955_),
    .ZN(_10071_));
 AND2_X1 _19381_ (.A1(_10070_),
    .A2(_10071_),
    .ZN(_10072_));
 NOR2_X1 _19382_ (.A1(_14835_),
    .A2(_09893_),
    .ZN(_10073_));
 CLKBUF_X3 _19383_ (.A(_10003_),
    .Z(_10074_));
 OAI21_X4 _19384_ (.A(_10013_),
    .B1(_09947_),
    .B2(_10074_),
    .ZN(_10075_));
 AOI21_X2 _19385_ (.A(_10073_),
    .B1(_10075_),
    .B2(_09949_),
    .ZN(_10076_));
 OAI221_X2 _19386_ (.A(_10067_),
    .B1(_10069_),
    .B2(_10072_),
    .C1(_10076_),
    .C2(_09830_),
    .ZN(_10077_));
 AND2_X2 _19387_ (.A1(_10066_),
    .A2(_10077_),
    .ZN(_10078_));
 NOR2_X2 _19388_ (.A1(_09890_),
    .A2(_09908_),
    .ZN(_10079_));
 OAI21_X1 _19389_ (.A(_09964_),
    .B1(_09831_),
    .B2(_10010_),
    .ZN(_10080_));
 NAND2_X1 _19390_ (.A1(_09951_),
    .A2(_10080_),
    .ZN(_10081_));
 OAI22_X1 _19391_ (.A1(_09928_),
    .A2(_09893_),
    .B1(_10030_),
    .B2(_10074_),
    .ZN(_10082_));
 AOI221_X2 _19392_ (.A(_10032_),
    .B1(_10079_),
    .B2(_10081_),
    .C1(_10082_),
    .C2(_09891_),
    .ZN(_10083_));
 NAND3_X1 _19393_ (.A1(_09940_),
    .A2(_09891_),
    .A3(_10023_),
    .ZN(_10084_));
 NAND2_X1 _19394_ (.A1(_09963_),
    .A2(_09924_),
    .ZN(_10085_));
 OAI21_X1 _19395_ (.A(_10084_),
    .B1(_10085_),
    .B2(net114),
    .ZN(_10086_));
 OAI22_X1 _19396_ (.A1(_10049_),
    .A2(_09904_),
    .B1(_09882_),
    .B2(_14835_),
    .ZN(_10087_));
 AOI22_X2 _19397_ (.A1(_14826_),
    .A2(_10086_),
    .B1(_10087_),
    .B2(net114),
    .ZN(_10088_));
 NOR2_X4 _19398_ (.A1(_14826_),
    .A2(_09948_),
    .ZN(_10089_));
 NOR2_X1 _19399_ (.A1(_09963_),
    .A2(_09951_),
    .ZN(_10090_));
 OAI21_X1 _19400_ (.A(_09951_),
    .B1(_09963_),
    .B2(net106),
    .ZN(_10091_));
 NAND2_X2 _19401_ (.A1(_09889_),
    .A2(_09851_),
    .ZN(_10092_));
 OAI21_X1 _19402_ (.A(_10091_),
    .B1(_10092_),
    .B2(_09928_),
    .ZN(_10093_));
 AOI221_X2 _19403_ (.A(_09984_),
    .B1(_10089_),
    .B2(_10090_),
    .C1(_10093_),
    .C2(_10025_),
    .ZN(_10094_));
 AOI21_X1 _19404_ (.A(_10083_),
    .B1(_10088_),
    .B2(_10094_),
    .ZN(_10095_));
 AOI221_X2 _19405_ (.A(_10036_),
    .B1(_10052_),
    .B2(_10078_),
    .C1(_10095_),
    .C2(_09806_),
    .ZN(_00041_));
 CLKBUF_X3 _19406_ (.A(_10023_),
    .Z(_10096_));
 NAND2_X1 _19407_ (.A1(_09863_),
    .A2(_09951_),
    .ZN(_10097_));
 OAI22_X1 _19408_ (.A1(_14856_),
    .A2(_10096_),
    .B1(_10097_),
    .B2(_10089_),
    .ZN(_10098_));
 NOR3_X2 _19409_ (.A1(net934),
    .A2(_14835_),
    .A3(_09949_),
    .ZN(_10099_));
 CLKBUF_X3 _19410_ (.A(_09938_),
    .Z(_10100_));
 MUX2_X1 _19411_ (.A(_14847_),
    .B(_10099_),
    .S(_10100_),
    .Z(_10101_));
 CLKBUF_X3 _19412_ (.A(_09996_),
    .Z(_10102_));
 NAND2_X1 _19413_ (.A1(_10102_),
    .A2(_10035_),
    .ZN(_10103_));
 OAI221_X1 _19414_ (.A(_09806_),
    .B1(_10019_),
    .B2(_10098_),
    .C1(_10101_),
    .C2(_10103_),
    .ZN(_10104_));
 NAND2_X1 _19415_ (.A1(net997),
    .A2(_10014_),
    .ZN(_10105_));
 AOI221_X1 _19416_ (.A(_09891_),
    .B1(_10029_),
    .B2(_09928_),
    .C1(_10105_),
    .C2(_10025_),
    .ZN(_10106_));
 NAND2_X1 _19417_ (.A1(_09894_),
    .A2(_09898_),
    .ZN(_10107_));
 NAND2_X4 _19418_ (.A1(_09854_),
    .A2(_09907_),
    .ZN(_10108_));
 OAI221_X1 _19419_ (.A(_10107_),
    .B1(_10108_),
    .B2(_09927_),
    .C1(_09933_),
    .C2(_10030_),
    .ZN(_10109_));
 CLKBUF_X3 _19420_ (.A(_09904_),
    .Z(_10110_));
 AOI21_X1 _19421_ (.A(_10106_),
    .B1(_10109_),
    .B2(_10110_),
    .ZN(_10111_));
 AOI21_X1 _19422_ (.A(_10104_),
    .B1(_10111_),
    .B2(_10033_),
    .ZN(_10112_));
 NAND4_X1 _19423_ (.A1(net114),
    .A2(_14851_),
    .A3(_09944_),
    .A4(_09947_),
    .ZN(_10113_));
 AOI211_X2 _19424_ (.A(_09984_),
    .B(_09903_),
    .C1(_09973_),
    .C2(_10010_),
    .ZN(_10114_));
 AOI21_X1 _19425_ (.A(_10037_),
    .B1(_10113_),
    .B2(_10114_),
    .ZN(_10115_));
 AOI21_X1 _19426_ (.A(_14844_),
    .B1(_09917_),
    .B2(net645),
    .ZN(_10116_));
 CLKBUF_X3 _19427_ (.A(_09932_),
    .Z(_10117_));
 OAI221_X1 _19428_ (.A(_09996_),
    .B1(_10117_),
    .B2(_09943_),
    .C1(_09977_),
    .C2(_09907_),
    .ZN(_10118_));
 OAI21_X2 _19429_ (.A(_10110_),
    .B1(_10116_),
    .B2(_10118_),
    .ZN(_10119_));
 NAND2_X1 _19430_ (.A1(_09854_),
    .A2(_09951_),
    .ZN(_10120_));
 AOI21_X1 _19431_ (.A(_09948_),
    .B1(_09932_),
    .B2(_09863_),
    .ZN(_10121_));
 NAND2_X1 _19432_ (.A1(_09917_),
    .A2(_09937_),
    .ZN(_10122_));
 AOI221_X2 _19433_ (.A(_09984_),
    .B1(_10120_),
    .B2(_10121_),
    .C1(_10122_),
    .C2(_09949_),
    .ZN(_10123_));
 AOI22_X1 _19434_ (.A1(_09907_),
    .A2(_14851_),
    .B1(_09905_),
    .B2(_09943_),
    .ZN(_10124_));
 OAI21_X1 _19435_ (.A(_10102_),
    .B1(_10100_),
    .B2(_10124_),
    .ZN(_10125_));
 OAI221_X2 _19436_ (.A(_10115_),
    .B1(_10119_),
    .B2(_10123_),
    .C1(_09967_),
    .C2(_10125_),
    .ZN(_10126_));
 AOI221_X1 _19437_ (.A(_09903_),
    .B1(_09914_),
    .B2(_09915_),
    .C1(_14826_),
    .C2(_10074_),
    .ZN(_10127_));
 AOI21_X1 _19438_ (.A(_10033_),
    .B1(_09965_),
    .B2(_10127_),
    .ZN(_10128_));
 OR3_X1 _19439_ (.A1(_14852_),
    .A2(_09904_),
    .A3(_10096_),
    .ZN(_10129_));
 AND2_X2 _19440_ (.A1(_09979_),
    .A2(_10014_),
    .ZN(_10130_));
 AOI21_X2 _19441_ (.A(_09894_),
    .B1(_09914_),
    .B2(_09915_),
    .ZN(_10131_));
 AOI21_X1 _19442_ (.A(_10131_),
    .B1(_10117_),
    .B2(_09943_),
    .ZN(_10132_));
 MUX2_X1 _19443_ (.A(_10130_),
    .B(_10132_),
    .S(_14844_),
    .Z(_10133_));
 OAI211_X2 _19444_ (.A(_10128_),
    .B(_10129_),
    .C1(_10035_),
    .C2(_10133_),
    .ZN(_10134_));
 NOR2_X1 _19445_ (.A1(_09984_),
    .A2(_09890_),
    .ZN(_10135_));
 AOI221_X2 _19446_ (.A(_09851_),
    .B1(_09905_),
    .B2(_09734_),
    .C1(_09989_),
    .C2(_09780_),
    .ZN(_10136_));
 AOI21_X1 _19447_ (.A(_10136_),
    .B1(_10117_),
    .B2(_14849_),
    .ZN(_10137_));
 NAND3_X1 _19448_ (.A1(_10074_),
    .A2(_10023_),
    .A3(_09992_),
    .ZN(_10138_));
 MUX2_X1 _19449_ (.A(_09948_),
    .B(_09897_),
    .S(_09863_),
    .Z(_10139_));
 OAI221_X2 _19450_ (.A(_10138_),
    .B1(_09965_),
    .B2(_10027_),
    .C1(net106),
    .C2(_10139_),
    .ZN(_10140_));
 AOI221_X2 _19451_ (.A(_09805_),
    .B1(_10137_),
    .B2(_10135_),
    .C1(_10140_),
    .C2(_10008_),
    .ZN(_10141_));
 AOI22_X2 _19452_ (.A1(_09931_),
    .A2(_10126_),
    .B1(_10134_),
    .B2(_10141_),
    .ZN(_10142_));
 OAI21_X4 _19453_ (.A(_09983_),
    .B1(_09948_),
    .B2(_09928_),
    .ZN(_10143_));
 AND2_X1 _19454_ (.A1(_10025_),
    .A2(_09980_),
    .ZN(_10144_));
 AOI21_X1 _19455_ (.A(_10143_),
    .B1(_10144_),
    .B2(_10097_),
    .ZN(_10145_));
 NOR3_X2 _19456_ (.A1(_10022_),
    .A2(_09887_),
    .A3(_09996_),
    .ZN(_10146_));
 OAI21_X1 _19457_ (.A(_09940_),
    .B1(_10023_),
    .B2(net619),
    .ZN(_10147_));
 NAND2_X1 _19458_ (.A1(_10032_),
    .A2(_09979_),
    .ZN(_10148_));
 OAI21_X1 _19459_ (.A(_09922_),
    .B1(_10147_),
    .B2(_10148_),
    .ZN(_10149_));
 NOR3_X1 _19460_ (.A1(_10145_),
    .A2(_10146_),
    .A3(_10149_),
    .ZN(_10150_));
 NAND2_X1 _19461_ (.A1(_09923_),
    .A2(_09959_),
    .ZN(_10151_));
 NAND2_X1 _19462_ (.A1(_09829_),
    .A2(_09890_),
    .ZN(_10152_));
 AOI21_X4 _19463_ (.A(net618),
    .B1(_09859_),
    .B2(_09861_),
    .ZN(_10153_));
 NOR3_X1 _19464_ (.A1(_10049_),
    .A2(_09887_),
    .A3(_10153_),
    .ZN(_10154_));
 NAND2_X1 _19465_ (.A1(_10010_),
    .A2(_09932_),
    .ZN(_10155_));
 AND3_X1 _19466_ (.A1(_09940_),
    .A2(_10097_),
    .A3(_10155_),
    .ZN(_10156_));
 NOR3_X1 _19467_ (.A1(_10152_),
    .A2(_10154_),
    .A3(_10156_),
    .ZN(_10157_));
 NAND3_X1 _19468_ (.A1(_14844_),
    .A2(_09917_),
    .A3(_09980_),
    .ZN(_10158_));
 NAND3_X1 _19469_ (.A1(_10049_),
    .A2(_10016_),
    .A3(net645),
    .ZN(_10159_));
 AOI21_X1 _19470_ (.A(_10019_),
    .B1(_10158_),
    .B2(_10159_),
    .ZN(_10160_));
 OR4_X1 _19471_ (.A1(_10150_),
    .A2(_10151_),
    .A3(_10157_),
    .A4(_10160_),
    .ZN(_10161_));
 AOI21_X2 _19472_ (.A(_10112_),
    .B1(_10142_),
    .B2(_10161_),
    .ZN(_00042_));
 NOR3_X4 _19473_ (.A1(net486),
    .A2(_09910_),
    .A3(_09911_),
    .ZN(_10162_));
 OAI21_X1 _19474_ (.A(_09784_),
    .B1(_10153_),
    .B2(_10162_),
    .ZN(_10163_));
 NAND3_X4 _19475_ (.A1(_10043_),
    .A2(_09944_),
    .A3(_09935_),
    .ZN(_10164_));
 AOI21_X4 _19476_ (.A(_09881_),
    .B1(_10164_),
    .B2(_10163_),
    .ZN(_10165_));
 OAI21_X1 _19477_ (.A(_09948_),
    .B1(_09897_),
    .B2(net112),
    .ZN(_10166_));
 AOI221_X2 _19478_ (.A(_09913_),
    .B1(_09898_),
    .B2(net112),
    .C1(_10166_),
    .C2(_09756_),
    .ZN(_10167_));
 AOI21_X4 _19479_ (.A(_10165_),
    .B1(_10167_),
    .B2(_09922_),
    .ZN(_10168_));
 NAND2_X1 _19480_ (.A1(_09884_),
    .A2(_09782_),
    .ZN(_10169_));
 NOR2_X2 _19481_ (.A1(_09781_),
    .A2(_10108_),
    .ZN(_10170_));
 NOR2_X1 _19482_ (.A1(_09924_),
    .A2(_10170_),
    .ZN(_10171_));
 AND2_X1 _19483_ (.A1(_10169_),
    .A2(_10171_),
    .ZN(_10172_));
 OR2_X2 _19484_ (.A1(_10064_),
    .A2(_10172_),
    .ZN(_10173_));
 NAND2_X1 _19485_ (.A1(_14842_),
    .A2(_14851_),
    .ZN(_10174_));
 NOR2_X1 _19486_ (.A1(_09955_),
    .A2(_10092_),
    .ZN(_10175_));
 AOI21_X1 _19487_ (.A(_09830_),
    .B1(_10174_),
    .B2(_10175_),
    .ZN(_10176_));
 AOI221_X2 _19488_ (.A(_10037_),
    .B1(_10168_),
    .B2(_10033_),
    .C1(_10173_),
    .C2(_10176_),
    .ZN(_10177_));
 OAI221_X1 _19489_ (.A(_09922_),
    .B1(_09927_),
    .B2(_09968_),
    .C1(_09893_),
    .C2(net110),
    .ZN(_10178_));
 OAI22_X1 _19490_ (.A1(_14844_),
    .A2(_09944_),
    .B1(_09992_),
    .B2(_10096_),
    .ZN(_10179_));
 AOI21_X1 _19491_ (.A(_10178_),
    .B1(_10179_),
    .B2(net114),
    .ZN(_10180_));
 NOR2_X1 _19492_ (.A1(_09959_),
    .A2(_09996_),
    .ZN(_10181_));
 BUF_X4 _19493_ (.A(_09891_),
    .Z(_10182_));
 OAI221_X1 _19494_ (.A(_10182_),
    .B1(_09893_),
    .B2(_09968_),
    .C1(_09944_),
    .C2(_14832_),
    .ZN(_10183_));
 AOI21_X1 _19495_ (.A(_14851_),
    .B1(_09917_),
    .B2(_09937_),
    .ZN(_10184_));
 OAI21_X1 _19496_ (.A(_10181_),
    .B1(_10183_),
    .B2(_10184_),
    .ZN(_10185_));
 OAI21_X1 _19497_ (.A(_14851_),
    .B1(_10110_),
    .B2(_14835_),
    .ZN(_10186_));
 AOI21_X1 _19498_ (.A(_10011_),
    .B1(_10100_),
    .B2(net619),
    .ZN(_10187_));
 AOI21_X1 _19499_ (.A(_10186_),
    .B1(_10187_),
    .B2(_10110_),
    .ZN(_10188_));
 NAND3_X1 _19500_ (.A1(net114),
    .A2(_10110_),
    .A3(_09973_),
    .ZN(_10189_));
 NOR2_X1 _19501_ (.A1(_09959_),
    .A2(_10033_),
    .ZN(_10190_));
 NOR3_X1 _19502_ (.A1(net113),
    .A2(_14835_),
    .A3(_09903_),
    .ZN(_10191_));
 NOR2_X1 _19503_ (.A1(_09935_),
    .A2(_09963_),
    .ZN(_10192_));
 AOI21_X1 _19504_ (.A(_09938_),
    .B1(_09903_),
    .B2(_10074_),
    .ZN(_10193_));
 AOI221_X2 _19505_ (.A(_10191_),
    .B1(_10192_),
    .B2(_10162_),
    .C1(_10193_),
    .C2(_10025_),
    .ZN(_10194_));
 NAND3_X1 _19506_ (.A1(_10189_),
    .A2(_10190_),
    .A3(_10194_),
    .ZN(_10195_));
 OAI221_X1 _19507_ (.A(_09923_),
    .B1(_10180_),
    .B2(_10185_),
    .C1(_10188_),
    .C2(_10195_),
    .ZN(_10196_));
 INV_X1 _19508_ (.A(_10181_),
    .ZN(_10197_));
 NOR3_X4 _19509_ (.A1(_09755_),
    .A2(_09846_),
    .A3(_09849_),
    .ZN(_10198_));
 NAND2_X1 _19510_ (.A1(_09940_),
    .A2(_10013_),
    .ZN(_10199_));
 MUX2_X1 _19511_ (.A(_09976_),
    .B(_09968_),
    .S(_09938_),
    .Z(_10200_));
 OAI221_X2 _19512_ (.A(_10182_),
    .B1(_10198_),
    .B2(_10199_),
    .C1(_10200_),
    .C2(_14851_),
    .ZN(_10201_));
 OAI21_X1 _19513_ (.A(_09937_),
    .B1(_10117_),
    .B2(_14842_),
    .ZN(_10202_));
 MUX2_X1 _19514_ (.A(_09907_),
    .B(net107),
    .S(_09932_),
    .Z(_10203_));
 MUX2_X1 _19515_ (.A(_10202_),
    .B(_10203_),
    .S(_10049_),
    .Z(_10204_));
 OAI21_X1 _19516_ (.A(_10201_),
    .B1(_10204_),
    .B2(_10110_),
    .ZN(_10205_));
 AOI21_X1 _19517_ (.A(_09955_),
    .B1(_09903_),
    .B2(_10074_),
    .ZN(_10206_));
 NOR2_X1 _19518_ (.A1(_10023_),
    .A2(_10206_),
    .ZN(_10207_));
 NOR3_X4 _19519_ (.A1(_09783_),
    .A2(_09876_),
    .A3(_09879_),
    .ZN(_10208_));
 NAND2_X1 _19520_ (.A1(_10074_),
    .A2(_10208_),
    .ZN(_10209_));
 MUX2_X1 _19521_ (.A(_09863_),
    .B(_09948_),
    .S(_09890_),
    .Z(_10210_));
 OAI21_X1 _19522_ (.A(_10209_),
    .B1(_10210_),
    .B2(_09900_),
    .ZN(_10211_));
 AOI21_X1 _19523_ (.A(_09924_),
    .B1(_09963_),
    .B2(_09989_),
    .ZN(_10212_));
 OAI22_X2 _19524_ (.A1(_14835_),
    .A2(_10085_),
    .B1(_10212_),
    .B2(_09940_),
    .ZN(_10213_));
 AOI221_X2 _19525_ (.A(_10207_),
    .B1(_10211_),
    .B2(_10096_),
    .C1(net114),
    .C2(_10213_),
    .ZN(_10214_));
 OAI21_X1 _19526_ (.A(_10190_),
    .B1(_09992_),
    .B2(_10035_),
    .ZN(_10215_));
 OAI221_X1 _19527_ (.A(_09931_),
    .B1(_10197_),
    .B2(_10205_),
    .C1(_10214_),
    .C2(_10215_),
    .ZN(_10216_));
 NOR2_X2 _19528_ (.A1(_10023_),
    .A2(_09992_),
    .ZN(_10217_));
 NOR2_X1 _19529_ (.A1(_09960_),
    .A2(_10217_),
    .ZN(_10218_));
 OAI21_X1 _19530_ (.A(_10218_),
    .B1(_09987_),
    .B2(_09884_),
    .ZN(_10219_));
 MUX2_X1 _19531_ (.A(_09900_),
    .B(_09756_),
    .S(_09831_),
    .Z(_10220_));
 NAND2_X1 _19532_ (.A1(_10010_),
    .A2(_09782_),
    .ZN(_10221_));
 AOI221_X1 _19533_ (.A(_10032_),
    .B1(_09938_),
    .B2(_10220_),
    .C1(_10221_),
    .C2(_10171_),
    .ZN(_10222_));
 OAI21_X1 _19534_ (.A(_09959_),
    .B1(_10110_),
    .B2(_10222_),
    .ZN(_10223_));
 NAND2_X1 _19535_ (.A1(_10074_),
    .A2(_09991_),
    .ZN(_10224_));
 NOR3_X1 _19536_ (.A1(_09894_),
    .A2(_09910_),
    .A3(_09911_),
    .ZN(_10225_));
 OAI21_X1 _19537_ (.A(_10049_),
    .B1(_10041_),
    .B2(_10225_),
    .ZN(_10226_));
 AOI21_X1 _19538_ (.A(_09830_),
    .B1(_10224_),
    .B2(_10226_),
    .ZN(_10227_));
 NAND2_X1 _19539_ (.A1(_09853_),
    .A2(_10096_),
    .ZN(_10228_));
 NAND3_X1 _19540_ (.A1(net106),
    .A2(_10032_),
    .A3(_10117_),
    .ZN(_10229_));
 AOI21_X1 _19541_ (.A(_14851_),
    .B1(_10228_),
    .B2(_10229_),
    .ZN(_10230_));
 OR2_X1 _19542_ (.A1(_10227_),
    .A2(_10230_),
    .ZN(_10231_));
 AOI22_X1 _19543_ (.A1(_10223_),
    .A2(_10219_),
    .B1(_10231_),
    .B2(_10110_),
    .ZN(_10232_));
 OAI22_X2 _19544_ (.A1(_10196_),
    .A2(_10177_),
    .B1(_10216_),
    .B2(_10232_),
    .ZN(_00043_));
 NAND2_X2 _19545_ (.A1(net997),
    .A2(_09935_),
    .ZN(_10233_));
 OAI221_X2 _19546_ (.A(_09904_),
    .B1(_10021_),
    .B2(_10233_),
    .C1(_10049_),
    .C2(net620),
    .ZN(_10234_));
 AOI21_X1 _19547_ (.A(_09924_),
    .B1(_14826_),
    .B2(net113),
    .ZN(_10235_));
 NAND2_X1 _19548_ (.A1(_09784_),
    .A2(_10043_),
    .ZN(_10236_));
 NOR2_X4 _19549_ (.A1(_10162_),
    .A2(_10153_),
    .ZN(_10237_));
 OAI221_X1 _19550_ (.A(_09881_),
    .B1(_10235_),
    .B2(_10236_),
    .C1(_10237_),
    .C2(_10025_),
    .ZN(_10238_));
 NAND4_X1 _19551_ (.A1(_10238_),
    .A2(_10234_),
    .A3(_10033_),
    .A4(_09806_),
    .ZN(_10239_));
 NAND2_X1 _19552_ (.A1(_09806_),
    .A2(_10102_),
    .ZN(_10240_));
 NAND2_X1 _19553_ (.A1(net112),
    .A2(_09862_),
    .ZN(_10241_));
 NOR3_X4 _19554_ (.A1(net647),
    .A2(_09910_),
    .A3(_09911_),
    .ZN(_10242_));
 NOR2_X4 _19555_ (.A1(_10242_),
    .A2(_09831_),
    .ZN(_10243_));
 OAI21_X4 _19556_ (.A(_10043_),
    .B1(_09852_),
    .B2(net689),
    .ZN(_10244_));
 AOI221_X2 _19557_ (.A(_09963_),
    .B1(_10243_),
    .B2(_10241_),
    .C1(_10244_),
    .C2(_09781_),
    .ZN(_10245_));
 NOR2_X1 _19558_ (.A1(net108),
    .A2(_09949_),
    .ZN(_10246_));
 NOR2_X1 _19559_ (.A1(net878),
    .A2(_09782_),
    .ZN(_10247_));
 OAI21_X1 _19560_ (.A(_10096_),
    .B1(_10246_),
    .B2(_10247_),
    .ZN(_10248_));
 AOI21_X2 _19561_ (.A(_10245_),
    .B1(_10248_),
    .B2(_10079_),
    .ZN(_10249_));
 OAI21_X2 _19562_ (.A(_10239_),
    .B1(_10240_),
    .B2(_10249_),
    .ZN(_10250_));
 AOI21_X1 _19563_ (.A(_09828_),
    .B1(_09914_),
    .B2(_09915_),
    .ZN(_10251_));
 AOI22_X2 _19564_ (.A1(_09736_),
    .A2(_09887_),
    .B1(_09955_),
    .B2(_10251_),
    .ZN(_10252_));
 AOI21_X1 _19565_ (.A(_10153_),
    .B1(_09938_),
    .B2(_09829_),
    .ZN(_10253_));
 AOI21_X1 _19566_ (.A(_09898_),
    .B1(_09973_),
    .B2(_10032_),
    .ZN(_10254_));
 OAI221_X2 _19567_ (.A(_10252_),
    .B1(_10253_),
    .B2(_10025_),
    .C1(_10254_),
    .C2(_09943_),
    .ZN(_10255_));
 AOI21_X1 _19568_ (.A(_09829_),
    .B1(_09862_),
    .B2(_09736_),
    .ZN(_10256_));
 AOI21_X1 _19569_ (.A(_10027_),
    .B1(_09924_),
    .B2(net878),
    .ZN(_10257_));
 OAI221_X2 _19570_ (.A(_10256_),
    .B1(_10257_),
    .B2(_09949_),
    .C1(_09853_),
    .C2(_09977_),
    .ZN(_10258_));
 INV_X1 _19571_ (.A(_14840_),
    .ZN(_10259_));
 MUX2_X1 _19572_ (.A(_10259_),
    .B(_09964_),
    .S(_09897_),
    .Z(_10260_));
 AOI21_X1 _19573_ (.A(_09891_),
    .B1(_10260_),
    .B2(_10032_),
    .ZN(_10261_));
 AOI22_X2 _19574_ (.A1(_10182_),
    .A2(_10255_),
    .B1(_10258_),
    .B2(_10261_),
    .ZN(_10262_));
 NAND2_X1 _19575_ (.A1(_09931_),
    .A2(_09959_),
    .ZN(_10263_));
 MUX2_X1 _19576_ (.A(_09965_),
    .B(_10070_),
    .S(_09889_),
    .Z(_10264_));
 OAI21_X1 _19577_ (.A(_09863_),
    .B1(_09756_),
    .B2(_10208_),
    .ZN(_10265_));
 AOI221_X2 _19578_ (.A(_09828_),
    .B1(_10264_),
    .B2(_09897_),
    .C1(_10265_),
    .C2(_10071_),
    .ZN(_10266_));
 NAND2_X1 _19579_ (.A1(_09828_),
    .A2(_09880_),
    .ZN(_10267_));
 NAND2_X1 _19580_ (.A1(net878),
    .A2(_09851_),
    .ZN(_10268_));
 AOI21_X4 _19581_ (.A(_09783_),
    .B1(_09886_),
    .B2(_09734_),
    .ZN(_10269_));
 AOI221_X2 _19582_ (.A(_10267_),
    .B1(_10268_),
    .B2(_10269_),
    .C1(_09948_),
    .C2(_09756_),
    .ZN(_10270_));
 MUX2_X1 _19583_ (.A(_09831_),
    .B(_09944_),
    .S(_09880_),
    .Z(_10271_));
 NOR3_X1 _19584_ (.A1(_09943_),
    .A2(_10032_),
    .A3(_10271_),
    .ZN(_10272_));
 OAI21_X1 _19585_ (.A(_09935_),
    .B1(_09924_),
    .B2(_09884_),
    .ZN(_10273_));
 AOI21_X1 _19586_ (.A(_10152_),
    .B1(_10273_),
    .B2(_10038_),
    .ZN(_10274_));
 NOR4_X2 _19587_ (.A1(_10274_),
    .A2(_10270_),
    .A3(_10272_),
    .A4(_10266_),
    .ZN(_10275_));
 NAND2_X2 _19588_ (.A1(_09923_),
    .A2(_10037_),
    .ZN(_10276_));
 OAI22_X2 _19589_ (.A1(_10262_),
    .A2(_10263_),
    .B1(_10275_),
    .B2(_10276_),
    .ZN(_10277_));
 AND2_X1 _19590_ (.A1(_09944_),
    .A2(_09937_),
    .ZN(_10278_));
 AOI221_X2 _19591_ (.A(_09984_),
    .B1(_10243_),
    .B2(_10039_),
    .C1(_10278_),
    .C2(_09782_),
    .ZN(_10279_));
 AOI221_X1 _19592_ (.A(_09829_),
    .B1(_09991_),
    .B2(_14826_),
    .C1(_10155_),
    .C2(_09782_),
    .ZN(_10280_));
 OAI21_X2 _19593_ (.A(_10035_),
    .B1(_10279_),
    .B2(_10280_),
    .ZN(_10281_));
 AOI21_X1 _19594_ (.A(_09781_),
    .B1(_10014_),
    .B2(_10016_),
    .ZN(_10282_));
 XNOR2_X1 _19595_ (.A(net107),
    .B(_09852_),
    .ZN(_10283_));
 AOI211_X2 _19596_ (.A(_09829_),
    .B(_10282_),
    .C1(_10283_),
    .C2(_09782_),
    .ZN(_10284_));
 AOI21_X1 _19597_ (.A(_10284_),
    .B1(_10040_),
    .B2(_10033_),
    .ZN(_10285_));
 OAI21_X2 _19598_ (.A(_10281_),
    .B1(_10285_),
    .B2(_10035_),
    .ZN(_10286_));
 INV_X1 _19599_ (.A(_10151_),
    .ZN(_10287_));
 AOI211_X2 _19600_ (.A(_10250_),
    .B(_10277_),
    .C1(_10286_),
    .C2(_10287_),
    .ZN(_00044_));
 NAND2_X1 _19601_ (.A1(_09931_),
    .A2(_09922_),
    .ZN(_10288_));
 NAND2_X1 _19602_ (.A1(_09943_),
    .A2(_10117_),
    .ZN(_10289_));
 OAI22_X1 _19603_ (.A1(_10289_),
    .A2(_10057_),
    .B1(_10108_),
    .B2(_09927_),
    .ZN(_10290_));
 AOI22_X1 _19604_ (.A1(_09928_),
    .A2(_09898_),
    .B1(_10221_),
    .B2(_10096_),
    .ZN(_10291_));
 NAND2_X1 _19605_ (.A1(_09931_),
    .A2(_10182_),
    .ZN(_10292_));
 OAI221_X1 _19606_ (.A(_09959_),
    .B1(_10288_),
    .B2(_10290_),
    .C1(_10291_),
    .C2(_10292_),
    .ZN(_10293_));
 NOR2_X2 _19607_ (.A1(net934),
    .A2(_09944_),
    .ZN(_10294_));
 OAI22_X1 _19608_ (.A1(_09999_),
    .A2(_10022_),
    .B1(_10147_),
    .B2(_10294_),
    .ZN(_10295_));
 AOI21_X1 _19609_ (.A(_10217_),
    .B1(_10289_),
    .B2(_14826_),
    .ZN(_10296_));
 MUX2_X1 _19610_ (.A(_10295_),
    .B(_10296_),
    .S(_10035_),
    .Z(_10297_));
 AOI21_X1 _19611_ (.A(_10293_),
    .B1(_10297_),
    .B2(_09923_),
    .ZN(_10298_));
 MUX2_X1 _19612_ (.A(_10010_),
    .B(_09736_),
    .S(_09932_),
    .Z(_10299_));
 AOI21_X1 _19613_ (.A(_09931_),
    .B1(_10208_),
    .B2(_10299_),
    .ZN(_10300_));
 OAI21_X1 _19614_ (.A(_10016_),
    .B1(_09893_),
    .B2(_09884_),
    .ZN(_10301_));
 OR3_X1 _19615_ (.A1(_09881_),
    .A2(_09888_),
    .A3(_10301_),
    .ZN(_10302_));
 NAND4_X1 _19616_ (.A1(_14844_),
    .A2(_09922_),
    .A3(_09916_),
    .A4(_10016_),
    .ZN(_10303_));
 AND3_X1 _19617_ (.A1(_10300_),
    .A2(_10302_),
    .A3(_10303_),
    .ZN(_10304_));
 NAND2_X1 _19618_ (.A1(_09890_),
    .A2(_09973_),
    .ZN(_10305_));
 AOI21_X1 _19619_ (.A(_09733_),
    .B1(_09880_),
    .B2(_09852_),
    .ZN(_10306_));
 AOI221_X1 _19620_ (.A(_14826_),
    .B1(_10305_),
    .B2(_10306_),
    .C1(_10092_),
    .C2(_10074_),
    .ZN(_10307_));
 NAND2_X1 _19621_ (.A1(_09881_),
    .A2(_10023_),
    .ZN(_10308_));
 AOI21_X1 _19622_ (.A(_09943_),
    .B1(_09977_),
    .B2(_10308_),
    .ZN(_10309_));
 AOI22_X1 _19623_ (.A1(_09894_),
    .A2(_10029_),
    .B1(_09991_),
    .B2(_14826_),
    .ZN(_10310_));
 NOR2_X1 _19624_ (.A1(_09922_),
    .A2(_10310_),
    .ZN(_10311_));
 NOR4_X1 _19625_ (.A1(_09923_),
    .A2(_10307_),
    .A3(_10309_),
    .A4(_10311_),
    .ZN(_10312_));
 NOR3_X2 _19626_ (.A1(_09959_),
    .A2(_10304_),
    .A3(_10312_),
    .ZN(_10313_));
 NAND2_X1 _19627_ (.A1(_09916_),
    .A2(_09979_),
    .ZN(_10314_));
 NAND2_X1 _19628_ (.A1(_09782_),
    .A2(_10314_),
    .ZN(_10315_));
 NAND3_X1 _19629_ (.A1(_09891_),
    .A2(_10224_),
    .A3(_10315_),
    .ZN(_10316_));
 OAI21_X1 _19630_ (.A(_10043_),
    .B1(_09851_),
    .B2(net878),
    .ZN(_10317_));
 AOI221_X2 _19631_ (.A(_09889_),
    .B1(_09989_),
    .B2(_09973_),
    .C1(_10317_),
    .C2(_09831_),
    .ZN(_10318_));
 NOR2_X1 _19632_ (.A1(_09795_),
    .A2(_10318_),
    .ZN(_10319_));
 NOR2_X1 _19633_ (.A1(_09782_),
    .A2(_10237_),
    .ZN(_10320_));
 OAI21_X1 _19634_ (.A(_09903_),
    .B1(_09935_),
    .B2(_09928_),
    .ZN(_10321_));
 OAI33_X1 _19635_ (.A1(_09904_),
    .A2(_09972_),
    .A3(_10320_),
    .B1(_10321_),
    .B2(_10294_),
    .B3(_09973_),
    .ZN(_10322_));
 AOI221_X2 _19636_ (.A(_09805_),
    .B1(_10319_),
    .B2(_10316_),
    .C1(_10322_),
    .C2(_09923_),
    .ZN(_10323_));
 OAI21_X1 _19637_ (.A(_09922_),
    .B1(_10100_),
    .B2(_09968_),
    .ZN(_10324_));
 AOI21_X1 _19638_ (.A(_10324_),
    .B1(_10062_),
    .B2(_10100_),
    .ZN(_10325_));
 OAI21_X1 _19639_ (.A(net645),
    .B1(_10117_),
    .B2(_09894_),
    .ZN(_10326_));
 NAND2_X1 _19640_ (.A1(_10049_),
    .A2(_10326_),
    .ZN(_10327_));
 NAND2_X1 _19641_ (.A1(_09937_),
    .A2(_10042_),
    .ZN(_10328_));
 AOI21_X1 _19642_ (.A(_10035_),
    .B1(_10327_),
    .B2(_10328_),
    .ZN(_10329_));
 NOR3_X1 _19643_ (.A1(_10263_),
    .A2(_10325_),
    .A3(_10329_),
    .ZN(_10330_));
 NOR2_X1 _19644_ (.A1(_10182_),
    .A2(_10217_),
    .ZN(_10331_));
 AOI21_X1 _19645_ (.A(_09881_),
    .B1(_09934_),
    .B2(_10025_),
    .ZN(_10332_));
 AOI22_X1 _19646_ (.A1(_09974_),
    .A2(_10331_),
    .B1(_10327_),
    .B2(_10332_),
    .ZN(_10333_));
 OAI21_X1 _19647_ (.A(_10102_),
    .B1(_10151_),
    .B2(_10333_),
    .ZN(_10334_));
 OAI33_X1 _19648_ (.A1(_10102_),
    .A2(_10298_),
    .A3(_10313_),
    .B1(_10323_),
    .B2(_10330_),
    .B3(_10334_),
    .ZN(_00045_));
 AOI21_X1 _19649_ (.A(_09783_),
    .B1(_09851_),
    .B2(_09884_),
    .ZN(_10335_));
 OAI21_X1 _19650_ (.A(_10043_),
    .B1(_09852_),
    .B2(_09854_),
    .ZN(_10336_));
 AOI221_X1 _19651_ (.A(_09828_),
    .B1(_10039_),
    .B2(_10335_),
    .C1(_10336_),
    .C2(_09784_),
    .ZN(_10337_));
 OAI221_X2 _19652_ (.A(_09933_),
    .B1(_09911_),
    .B2(_09910_),
    .C1(_09863_),
    .C2(_09781_),
    .ZN(_10338_));
 OR3_X1 _19653_ (.A1(_14845_),
    .A2(_14854_),
    .A3(_09897_),
    .ZN(_10339_));
 AOI21_X1 _19654_ (.A(_09996_),
    .B1(_10338_),
    .B2(_10339_),
    .ZN(_10340_));
 NOR3_X1 _19655_ (.A1(_10182_),
    .A2(_10337_),
    .A3(_10340_),
    .ZN(_10341_));
 OAI21_X1 _19656_ (.A(_10014_),
    .B1(_09852_),
    .B2(_09884_),
    .ZN(_10342_));
 NAND2_X1 _19657_ (.A1(_09948_),
    .A2(_10342_),
    .ZN(_10343_));
 AOI21_X1 _19658_ (.A(_09983_),
    .B1(_10029_),
    .B2(_09853_),
    .ZN(_10344_));
 OR2_X2 _19659_ (.A1(_10153_),
    .A2(_10198_),
    .ZN(_10345_));
 OAI21_X1 _19660_ (.A(_09937_),
    .B1(_10108_),
    .B2(_09851_),
    .ZN(_10346_));
 MUX2_X1 _19661_ (.A(_10345_),
    .B(_10346_),
    .S(_09831_),
    .Z(_10347_));
 AOI221_X2 _19662_ (.A(_09963_),
    .B1(_10343_),
    .B2(_10344_),
    .C1(_10347_),
    .C2(_09984_),
    .ZN(_10348_));
 NOR3_X1 _19663_ (.A1(_10348_),
    .A2(_10341_),
    .A3(_10276_),
    .ZN(_10349_));
 OAI21_X1 _19664_ (.A(_09890_),
    .B1(_10198_),
    .B2(net107),
    .ZN(_10350_));
 AOI21_X1 _19665_ (.A(_09948_),
    .B1(_09880_),
    .B2(_09862_),
    .ZN(_10351_));
 OAI22_X2 _19666_ (.A1(_14835_),
    .A2(_10092_),
    .B1(_10237_),
    .B2(_09890_),
    .ZN(_10352_));
 AOI221_X2 _19667_ (.A(_09829_),
    .B1(_10350_),
    .B2(_10351_),
    .C1(_10352_),
    .C2(_09949_),
    .ZN(_10353_));
 NOR2_X1 _19668_ (.A1(_09992_),
    .A2(_10308_),
    .ZN(_10354_));
 AOI21_X1 _19669_ (.A(_10089_),
    .B1(_09862_),
    .B2(net108),
    .ZN(_10355_));
 AOI21_X1 _19670_ (.A(_10198_),
    .B1(_09905_),
    .B2(_10074_),
    .ZN(_10356_));
 OAI21_X1 _19671_ (.A(_10355_),
    .B1(_10356_),
    .B2(_14842_),
    .ZN(_10357_));
 AOI21_X1 _19672_ (.A(_10354_),
    .B1(_10357_),
    .B2(_10182_),
    .ZN(_10358_));
 OAI22_X1 _19673_ (.A1(_09904_),
    .A2(_10089_),
    .B1(_10155_),
    .B2(_09940_),
    .ZN(_10359_));
 AOI21_X1 _19674_ (.A(_09996_),
    .B1(_10359_),
    .B2(_14832_),
    .ZN(_10360_));
 AOI21_X1 _19675_ (.A(_10353_),
    .B1(_10358_),
    .B2(_10360_),
    .ZN(_10361_));
 NOR2_X1 _19676_ (.A1(_10198_),
    .A2(_10011_),
    .ZN(_10362_));
 OAI221_X1 _19677_ (.A(_10008_),
    .B1(_10362_),
    .B2(_14844_),
    .C1(_09927_),
    .C2(net110),
    .ZN(_10363_));
 NOR2_X1 _19678_ (.A1(_09829_),
    .A2(_09963_),
    .ZN(_10364_));
 AOI21_X1 _19679_ (.A(_10153_),
    .B1(_10117_),
    .B2(_09894_),
    .ZN(_10365_));
 OAI22_X1 _19680_ (.A1(net114),
    .A2(_09927_),
    .B1(_10365_),
    .B2(_14844_),
    .ZN(_10366_));
 AOI21_X1 _19681_ (.A(_10143_),
    .B1(_09905_),
    .B2(net113),
    .ZN(_10367_));
 NOR2_X1 _19682_ (.A1(_14846_),
    .A2(_09984_),
    .ZN(_10368_));
 NOR2_X1 _19683_ (.A1(_09884_),
    .A2(_09784_),
    .ZN(_10369_));
 NAND2_X1 _19684_ (.A1(_09829_),
    .A2(_09924_),
    .ZN(_10370_));
 NOR2_X1 _19685_ (.A1(net107),
    .A2(_09781_),
    .ZN(_10371_));
 OAI33_X1 _19686_ (.A1(_10367_),
    .A2(_10100_),
    .A3(_10368_),
    .B1(_10369_),
    .B2(_10370_),
    .B3(_10371_),
    .ZN(_10372_));
 AOI22_X1 _19687_ (.A1(_10364_),
    .A2(_10366_),
    .B1(_10035_),
    .B2(_10372_),
    .ZN(_10373_));
 NAND3_X1 _19688_ (.A1(_10373_),
    .A2(_10363_),
    .A3(_09959_),
    .ZN(_10374_));
 OAI21_X1 _19689_ (.A(_10117_),
    .B1(_09940_),
    .B2(net110),
    .ZN(_10375_));
 OAI221_X2 _19690_ (.A(_10008_),
    .B1(_10099_),
    .B2(_10375_),
    .C1(_10100_),
    .C2(_14847_),
    .ZN(_10376_));
 OAI21_X1 _19691_ (.A(_09784_),
    .B1(_09951_),
    .B2(_10108_),
    .ZN(_10377_));
 OAI221_X1 _19692_ (.A(_09975_),
    .B1(_10122_),
    .B2(_09949_),
    .C1(_10377_),
    .C2(_10294_),
    .ZN(_10378_));
 NOR2_X1 _19693_ (.A1(net934),
    .A2(_09955_),
    .ZN(_10379_));
 OAI221_X1 _19694_ (.A(_10364_),
    .B1(_10379_),
    .B2(_09938_),
    .C1(_09893_),
    .C2(_09894_),
    .ZN(_10380_));
 NAND2_X1 _19695_ (.A1(_09781_),
    .A2(_10038_),
    .ZN(_10381_));
 OAI21_X1 _19696_ (.A(_09937_),
    .B1(_09924_),
    .B2(_09863_),
    .ZN(_10382_));
 OAI221_X1 _19697_ (.A(_10135_),
    .B1(_10381_),
    .B2(_10294_),
    .C1(_10382_),
    .C2(_09940_),
    .ZN(_10383_));
 AND4_X2 _19698_ (.A1(_10037_),
    .A2(_10378_),
    .A3(_10380_),
    .A4(_10383_),
    .ZN(_10384_));
 AOI21_X2 _19699_ (.A(_09923_),
    .B1(_10376_),
    .B2(_10384_),
    .ZN(_10385_));
 AOI221_X1 _19700_ (.A(_10349_),
    .B1(_10361_),
    .B2(_10287_),
    .C1(_10374_),
    .C2(_10385_),
    .ZN(_00046_));
 NAND3_X1 _19701_ (.A1(_09853_),
    .A2(_10049_),
    .A3(_10100_),
    .ZN(_10386_));
 OAI21_X1 _19702_ (.A(_10386_),
    .B1(_10100_),
    .B2(_14840_),
    .ZN(_10387_));
 OAI21_X1 _19703_ (.A(_10110_),
    .B1(_10096_),
    .B2(_10379_),
    .ZN(_10388_));
 OAI221_X1 _19704_ (.A(_09806_),
    .B1(_10267_),
    .B2(_10387_),
    .C1(_10388_),
    .C2(_10069_),
    .ZN(_10389_));
 OAI21_X1 _19705_ (.A(_10117_),
    .B1(_09940_),
    .B2(_09884_),
    .ZN(_10390_));
 OAI221_X1 _19706_ (.A(_09922_),
    .B1(_10002_),
    .B2(_10390_),
    .C1(_10100_),
    .C2(_14854_),
    .ZN(_10391_));
 OAI211_X2 _19707_ (.A(_10025_),
    .B(_10013_),
    .C1(_10023_),
    .C2(net108),
    .ZN(_10392_));
 NAND3_X1 _19708_ (.A1(_10182_),
    .A2(_10047_),
    .A3(_10392_),
    .ZN(_10393_));
 AND3_X1 _19709_ (.A1(_10102_),
    .A2(_10391_),
    .A3(_10393_),
    .ZN(_10394_));
 OR2_X1 _19710_ (.A1(_10389_),
    .A2(_10394_),
    .ZN(_10395_));
 NOR2_X1 _19711_ (.A1(_09923_),
    .A2(_10033_),
    .ZN(_10396_));
 AOI21_X1 _19712_ (.A(_09898_),
    .B1(_10096_),
    .B2(_09881_),
    .ZN(_10397_));
 NOR3_X1 _19713_ (.A1(net108),
    .A2(_14826_),
    .A3(_10397_),
    .ZN(_10398_));
 NAND4_X1 _19714_ (.A1(_09943_),
    .A2(_09891_),
    .A3(_10023_),
    .A4(_09905_),
    .ZN(_10399_));
 OAI221_X1 _19715_ (.A(_10399_),
    .B1(_09904_),
    .B2(_14844_),
    .C1(net106),
    .C2(_09977_),
    .ZN(_10400_));
 OAI21_X1 _19716_ (.A(_10396_),
    .B1(_10398_),
    .B2(_10400_),
    .ZN(_10401_));
 NAND2_X1 _19717_ (.A1(_09931_),
    .A2(_10033_),
    .ZN(_10402_));
 OAI21_X1 _19718_ (.A(_09947_),
    .B1(_09927_),
    .B2(_14835_),
    .ZN(_10403_));
 NAND2_X1 _19719_ (.A1(_10182_),
    .A2(_10403_),
    .ZN(_10404_));
 AOI21_X1 _19720_ (.A(_09736_),
    .B1(_09917_),
    .B2(_09893_),
    .ZN(_10405_));
 AOI21_X1 _19721_ (.A(_10405_),
    .B1(_09887_),
    .B2(_09943_),
    .ZN(_10406_));
 NOR2_X1 _19722_ (.A1(_10029_),
    .A2(_10217_),
    .ZN(_10407_));
 OAI221_X1 _19723_ (.A(_10404_),
    .B1(_10406_),
    .B2(_10182_),
    .C1(net108),
    .C2(_10407_),
    .ZN(_10408_));
 OAI22_X4 _19724_ (.A1(net619),
    .A2(_09882_),
    .B1(_10244_),
    .B2(_14851_),
    .ZN(_10409_));
 OAI21_X4 _19725_ (.A(_10067_),
    .B1(_10409_),
    .B2(_10102_),
    .ZN(_10410_));
 AND2_X1 _19726_ (.A1(_09917_),
    .A2(net645),
    .ZN(_10411_));
 AOI221_X2 _19727_ (.A(_09830_),
    .B1(_09980_),
    .B2(_10269_),
    .C1(_10411_),
    .C2(_14844_),
    .ZN(_10412_));
 OAI221_X2 _19728_ (.A(_10401_),
    .B1(_10402_),
    .B2(_10408_),
    .C1(_10410_),
    .C2(_10412_),
    .ZN(_10413_));
 AOI21_X1 _19729_ (.A(_09887_),
    .B1(_10089_),
    .B2(_10096_),
    .ZN(_10414_));
 OAI221_X1 _19730_ (.A(_09830_),
    .B1(_09927_),
    .B2(_09976_),
    .C1(_10414_),
    .C2(net108),
    .ZN(_10415_));
 OAI221_X1 _19731_ (.A(_09996_),
    .B1(_09927_),
    .B2(_14842_),
    .C1(_10030_),
    .C2(net110),
    .ZN(_10416_));
 AOI21_X1 _19732_ (.A(_10073_),
    .B1(_10415_),
    .B2(_10416_),
    .ZN(_10417_));
 OAI21_X1 _19733_ (.A(_09959_),
    .B1(_10046_),
    .B2(_10417_),
    .ZN(_10418_));
 NOR2_X1 _19734_ (.A1(_10033_),
    .A2(_10242_),
    .ZN(_10419_));
 AOI21_X1 _19735_ (.A(_10035_),
    .B1(_10338_),
    .B2(_10419_),
    .ZN(_10420_));
 NOR2_X1 _19736_ (.A1(_10198_),
    .A2(_10153_),
    .ZN(_10421_));
 AOI221_X1 _19737_ (.A(_09999_),
    .B1(_10108_),
    .B2(_09973_),
    .C1(_10421_),
    .C2(_10049_),
    .ZN(_10422_));
 OAI21_X1 _19738_ (.A(_10420_),
    .B1(_10422_),
    .B2(_10102_),
    .ZN(_10423_));
 OAI21_X1 _19739_ (.A(_14851_),
    .B1(_10131_),
    .B2(_09934_),
    .ZN(_10424_));
 NOR2_X1 _19740_ (.A1(_10102_),
    .A2(_10015_),
    .ZN(_10425_));
 AOI21_X1 _19741_ (.A(_10247_),
    .B1(_10269_),
    .B2(_10038_),
    .ZN(_10426_));
 AOI22_X1 _19742_ (.A1(_10424_),
    .A2(_10425_),
    .B1(_10426_),
    .B2(_10102_),
    .ZN(_10427_));
 OAI21_X1 _19743_ (.A(_10423_),
    .B1(_10427_),
    .B2(_10110_),
    .ZN(_10428_));
 OAI221_X1 _19744_ (.A(_10395_),
    .B1(_10413_),
    .B2(_10418_),
    .C1(_10428_),
    .C2(_10276_),
    .ZN(_00047_));
 INV_X1 _19745_ (.A(net796),
    .ZN(_10429_));
 NOR2_X1 _19746_ (.A1(_10429_),
    .A2(net610),
    .ZN(_10430_));
 NOR2_X1 _19747_ (.A1(net797),
    .A2(_09728_),
    .ZN(_10431_));
 BUF_X4 _19748_ (.A(\sa02_sr[7] ),
    .Z(_10432_));
 BUF_X1 rebuffer53 (.A(_15167_),
    .Z(net537));
 XOR2_X2 _19750_ (.A(\sa12_sr[7] ),
    .B(_10432_),
    .Z(_10434_));
 BUF_X4 clone95 (.A(_04987_),
    .Z(net95));
 BUF_X8 clone96 (.A(net1153),
    .Z(net96));
 XNOR2_X2 _19753_ (.A(\sa12_sr[1] ),
    .B(\sa20_sub[1] ),
    .ZN(_10437_));
 XNOR2_X1 _19754_ (.A(_10434_),
    .B(_10437_),
    .ZN(_10438_));
 BUF_X4 _19755_ (.A(\sa02_sr[0] ),
    .Z(_10439_));
 BUF_X4 clone5 (.A(net1233),
    .Z(net5));
 BUF_X4 clone153 (.A(net512),
    .Z(net153));
 XOR2_X2 _19758_ (.A(net595),
    .B(net531),
    .Z(_10442_));
 XNOR2_X2 _19759_ (.A(_10439_),
    .B(_10442_),
    .ZN(_10443_));
 XNOR2_X2 _19760_ (.A(_10438_),
    .B(_10443_),
    .ZN(_10444_));
 MUX2_X2 _19761_ (.A(_10430_),
    .B(_10431_),
    .S(_10444_),
    .Z(_10445_));
 NOR3_X2 _19762_ (.A1(net796),
    .A2(_09100_),
    .A3(_00446_),
    .ZN(_10446_));
 NOR2_X1 _19763_ (.A1(_10429_),
    .A2(_09075_),
    .ZN(_10447_));
 AOI21_X4 _19764_ (.A(_10446_),
    .B1(_10447_),
    .B2(_00446_),
    .ZN(_10448_));
 INV_X2 _19765_ (.A(_10448_),
    .ZN(_10449_));
 NOR2_X4 _19766_ (.A1(_10445_),
    .A2(_10449_),
    .ZN(_10450_));
 INV_X1 _19767_ (.A(_10450_),
    .ZN(_10451_));
 BUF_X4 _19768_ (.A(_10451_),
    .Z(_10452_));
 BUF_X8 _19769_ (.A(_10452_),
    .Z(_14864_));
 BUF_X4 _19770_ (.A(\sa31_sub[0] ),
    .Z(_10453_));
 BUF_X4 clone57 (.A(net792),
    .Z(net57));
 XNOR2_X2 _19772_ (.A(net598),
    .B(\sa12_sr[0] ),
    .ZN(_10455_));
 XNOR2_X1 _19773_ (.A(_10453_),
    .B(net573),
    .ZN(_10456_));
 NAND3_X1 _19774_ (.A1(net793),
    .A2(_09023_),
    .A3(_10434_),
    .ZN(_10457_));
 XNOR2_X2 _19775_ (.A(_10432_),
    .B(net549),
    .ZN(_10458_));
 NOR2_X1 _19776_ (.A1(net793),
    .A2(_09027_),
    .ZN(_10459_));
 NAND2_X1 _19777_ (.A1(_10458_),
    .A2(_10459_),
    .ZN(_10460_));
 AOI21_X1 _19778_ (.A(_10456_),
    .B1(_10457_),
    .B2(_10460_),
    .ZN(_10461_));
 XOR2_X1 _19779_ (.A(_10453_),
    .B(net573),
    .Z(_10462_));
 NAND2_X1 _19780_ (.A1(_10434_),
    .A2(_10459_),
    .ZN(_10463_));
 NAND3_X1 _19781_ (.A1(net793),
    .A2(_09194_),
    .A3(_10458_),
    .ZN(_10464_));
 AOI21_X1 _19782_ (.A(_10462_),
    .B1(_10463_),
    .B2(_10464_),
    .ZN(_10465_));
 INV_X1 _19783_ (.A(net793),
    .ZN(_10466_));
 NAND3_X1 _19784_ (.A1(_10466_),
    .A2(_09727_),
    .A3(_00447_),
    .ZN(_10467_));
 NAND2_X1 _19785_ (.A1(net793),
    .A2(_09028_),
    .ZN(_10468_));
 OAI21_X1 _19786_ (.A(_10467_),
    .B1(_10468_),
    .B2(_00447_),
    .ZN(_10469_));
 OR3_X1 _19787_ (.A1(_10461_),
    .A2(_10465_),
    .A3(_10469_),
    .ZN(_10470_));
 BUF_X4 _19788_ (.A(_10470_),
    .Z(_10471_));
 INV_X2 _19789_ (.A(_10471_),
    .ZN(_10472_));
 BUF_X8 _19790_ (.A(_10472_),
    .Z(_10473_));
 BUF_X4 _19791_ (.A(_10473_),
    .Z(_14867_));
 BUF_X4 clone133 (.A(net174),
    .Z(net133));
 BUF_X4 _19793_ (.A(\sa31_sub[2] ),
    .Z(_10475_));
 XOR2_X2 _19794_ (.A(net533),
    .B(_10475_),
    .Z(_10476_));
 XOR2_X1 _19795_ (.A(net585),
    .B(_10476_),
    .Z(_10477_));
 BUF_X4 _19796_ (.A(\sa12_sr[2] ),
    .Z(_10478_));
 BUF_X4 _19797_ (.A(\sa20_sub[2] ),
    .Z(_10479_));
 XOR2_X2 _19798_ (.A(_10478_),
    .B(_10479_),
    .Z(_10480_));
 NAND3_X1 _19799_ (.A1(_06637_),
    .A2(_09011_),
    .A3(_10480_),
    .ZN(_10481_));
 XNOR2_X2 _19800_ (.A(_10478_),
    .B(_10479_),
    .ZN(_10482_));
 NOR2_X1 _19801_ (.A1(_06637_),
    .A2(_08992_),
    .ZN(_10483_));
 NAND2_X1 _19802_ (.A1(_10482_),
    .A2(_10483_),
    .ZN(_10484_));
 AOI21_X2 _19803_ (.A(_10477_),
    .B1(_10481_),
    .B2(_10484_),
    .ZN(_10485_));
 XNOR2_X1 _19804_ (.A(net585),
    .B(_10476_),
    .ZN(_10486_));
 NAND2_X1 _19805_ (.A1(_10480_),
    .A2(_10483_),
    .ZN(_10487_));
 NAND3_X1 _19806_ (.A1(_06637_),
    .A2(_09022_),
    .A3(_10482_),
    .ZN(_10488_));
 AOI21_X2 _19807_ (.A(_10486_),
    .B1(_10487_),
    .B2(_10488_),
    .ZN(_10489_));
 INV_X1 _19808_ (.A(_06637_),
    .ZN(_10490_));
 NAND3_X1 _19809_ (.A1(_10490_),
    .A2(_09027_),
    .A3(_00448_),
    .ZN(_10491_));
 NAND2_X1 _19810_ (.A1(_06637_),
    .A2(_09027_),
    .ZN(_10492_));
 OAI21_X2 _19811_ (.A(_10491_),
    .B1(_10492_),
    .B2(_00448_),
    .ZN(_10493_));
 NOR3_X4 _19812_ (.A1(_10485_),
    .A2(_10489_),
    .A3(_10493_),
    .ZN(_10494_));
 INV_X4 _19813_ (.A(_10494_),
    .ZN(_10495_));
 BUF_X4 _19814_ (.A(_10495_),
    .Z(_10496_));
 BUF_X4 _19815_ (.A(_10496_),
    .Z(_10497_));
 BUF_X4 _19816_ (.A(_10497_),
    .Z(_10498_));
 BUF_X4 _19817_ (.A(_10498_),
    .Z(_10499_));
 BUF_X4 _19818_ (.A(_10499_),
    .Z(_14883_));
 BUF_X4 _19819_ (.A(_10471_),
    .Z(_14858_));
 BUF_X4 _19820_ (.A(_10494_),
    .Z(_10500_));
 BUF_X4 _19821_ (.A(_10500_),
    .Z(_10501_));
 BUF_X4 _19822_ (.A(_10501_),
    .Z(_14876_));
 CLKBUF_X3 _19823_ (.A(\sa12_sr[6] ),
    .Z(_10502_));
 BUF_X4 _19824_ (.A(\sa20_sub[7] ),
    .Z(_10503_));
 XNOR2_X2 _19825_ (.A(\sa12_sr[7] ),
    .B(_10503_),
    .ZN(_10504_));
 BUF_X2 _19826_ (.A(\sa02_sr[6] ),
    .Z(_10505_));
 BUF_X8 _19827_ (.A(\sa31_sub[7] ),
    .Z(_10506_));
 XNOR2_X1 _19828_ (.A(_10505_),
    .B(net712),
    .ZN(_10507_));
 XNOR2_X1 _19829_ (.A(_10504_),
    .B(_10507_),
    .ZN(_10508_));
 XNOR2_X1 _19830_ (.A(_10502_),
    .B(_10508_),
    .ZN(_10509_));
 MUX2_X2 _19831_ (.A(\text_in_r[63] ),
    .B(_10509_),
    .S(_09158_),
    .Z(_10510_));
 XOR2_X2 _19832_ (.A(_06710_),
    .B(_10510_),
    .Z(_10511_));
 CLKBUF_X3 _19833_ (.A(\sa31_sub[6] ),
    .Z(_10512_));
 BUF_X2 _19834_ (.A(\sa20_sub[6] ),
    .Z(_10513_));
 XNOR2_X2 _19835_ (.A(_10502_),
    .B(_10513_),
    .ZN(_10514_));
 BUF_X4 _19836_ (.A(\sa12_sr[5] ),
    .Z(_10515_));
 BUF_X2 _19837_ (.A(\sa02_sr[5] ),
    .Z(_10516_));
 XNOR2_X2 _19838_ (.A(_10515_),
    .B(_10516_),
    .ZN(_10517_));
 XNOR2_X1 _19839_ (.A(_10514_),
    .B(_10517_),
    .ZN(_10518_));
 XNOR2_X1 _19840_ (.A(_10512_),
    .B(_10518_),
    .ZN(_10519_));
 MUX2_X2 _19841_ (.A(\text_in_r[62] ),
    .B(_10519_),
    .S(_09195_),
    .Z(_10520_));
 XNOR2_X2 _19842_ (.A(_06696_),
    .B(_10520_),
    .ZN(_10521_));
 NAND2_X2 _19843_ (.A1(_10511_),
    .A2(_10521_),
    .ZN(_10522_));
 BUF_X2 _19844_ (.A(\sa20_sub[5] ),
    .Z(_10523_));
 CLKBUF_X3 _19845_ (.A(\sa31_sub[5] ),
    .Z(_10524_));
 XNOR2_X2 _19846_ (.A(_10523_),
    .B(_10524_),
    .ZN(_10525_));
 CLKBUF_X3 _19847_ (.A(\sa12_sr[4] ),
    .Z(_10526_));
 BUF_X2 _19848_ (.A(\sa02_sr[4] ),
    .Z(_10527_));
 XNOR2_X2 _19849_ (.A(_10526_),
    .B(_10527_),
    .ZN(_10528_));
 XNOR2_X1 _19850_ (.A(_10525_),
    .B(_10528_),
    .ZN(_10529_));
 XNOR2_X1 _19851_ (.A(_10515_),
    .B(_10529_),
    .ZN(_10530_));
 MUX2_X2 _19852_ (.A(\text_in_r[61] ),
    .B(_10530_),
    .S(_09076_),
    .Z(_10531_));
 XOR2_X2 _19853_ (.A(_06687_),
    .B(_10531_),
    .Z(_10532_));
 BUF_X4 _19854_ (.A(_10532_),
    .Z(_10533_));
 BUF_X4 _19855_ (.A(_10533_),
    .Z(_10534_));
 BUF_X2 _19856_ (.A(\sa02_sr[3] ),
    .Z(_10535_));
 BUF_X2 _19857_ (.A(\sa20_sub[4] ),
    .Z(_10536_));
 XNOR2_X2 _19858_ (.A(_10535_),
    .B(_10536_),
    .ZN(_10537_));
 XNOR2_X2 _19859_ (.A(_10432_),
    .B(_10537_),
    .ZN(_10538_));
 BUF_X2 _19860_ (.A(\sa12_sr[3] ),
    .Z(_10539_));
 XOR2_X2 _19861_ (.A(net552),
    .B(_10539_),
    .Z(_10540_));
 CLKBUF_X3 _19862_ (.A(\sa31_sub[4] ),
    .Z(_10541_));
 XOR2_X1 _19863_ (.A(_10526_),
    .B(_10541_),
    .Z(_10542_));
 XNOR2_X1 _19864_ (.A(_10540_),
    .B(_10542_),
    .ZN(_10543_));
 XNOR2_X1 _19865_ (.A(_10538_),
    .B(_10543_),
    .ZN(_10544_));
 MUX2_X2 _19866_ (.A(\text_in_r[60] ),
    .B(_10544_),
    .S(_09075_),
    .Z(_10545_));
 XOR2_X2 _19867_ (.A(_06672_),
    .B(_10545_),
    .Z(_10546_));
 INV_X1 _19868_ (.A(_06656_),
    .ZN(_10547_));
 NAND2_X1 _19869_ (.A1(_10547_),
    .A2(_09076_),
    .ZN(_10548_));
 NAND2_X1 _19870_ (.A1(_06656_),
    .A2(_09076_),
    .ZN(_10549_));
 BUF_X4 _19871_ (.A(\sa02_sr[2] ),
    .Z(_10550_));
 BUF_X2 _19872_ (.A(\sa20_sub[3] ),
    .Z(_10551_));
 XNOR2_X1 _19873_ (.A(_10550_),
    .B(_10551_),
    .ZN(_10552_));
 XNOR2_X2 _19874_ (.A(_10432_),
    .B(_10552_),
    .ZN(_10553_));
 BUF_X4 _19875_ (.A(\sa31_sub[3] ),
    .Z(_10554_));
 XNOR2_X1 _19876_ (.A(_10478_),
    .B(_10554_),
    .ZN(_10555_));
 XNOR2_X1 _19877_ (.A(_10540_),
    .B(_10555_),
    .ZN(_10556_));
 XNOR2_X2 _19878_ (.A(_10553_),
    .B(_10556_),
    .ZN(_10557_));
 MUX2_X2 _19879_ (.A(_10548_),
    .B(_10549_),
    .S(_10557_),
    .Z(_10558_));
 OR3_X2 _19880_ (.A1(_10547_),
    .A2(net949),
    .A3(\text_in_r[59] ),
    .ZN(_10559_));
 NAND3_X2 _19881_ (.A1(_10547_),
    .A2(net610),
    .A3(\text_in_r[59] ),
    .ZN(_10560_));
 AND2_X1 _19882_ (.A1(_10559_),
    .A2(_10560_),
    .ZN(_10561_));
 BUF_X4 _19883_ (.A(_10561_),
    .Z(_10562_));
 AOI21_X4 _19884_ (.A(_10494_),
    .B1(_10558_),
    .B2(_10562_),
    .ZN(_10563_));
 BUF_X4 _19885_ (.A(_14870_),
    .Z(_10564_));
 NOR2_X1 _19886_ (.A1(_06656_),
    .A2(_09028_),
    .ZN(_10565_));
 NOR2_X1 _19887_ (.A1(_10547_),
    .A2(_09028_),
    .ZN(_10566_));
 MUX2_X1 _19888_ (.A(_10565_),
    .B(_10566_),
    .S(_10557_),
    .Z(_10567_));
 BUF_X4 _19889_ (.A(_10567_),
    .Z(_10568_));
 NAND2_X4 _19890_ (.A1(_10559_),
    .A2(_10560_),
    .ZN(_10569_));
 NOR3_X4 _19891_ (.A1(net599),
    .A2(_10568_),
    .A3(_10569_),
    .ZN(_10570_));
 BUF_X4 _19892_ (.A(_09118_),
    .Z(_10571_));
 NAND2_X1 _19893_ (.A1(net797),
    .A2(_10571_),
    .ZN(_10572_));
 NAND2_X1 _19894_ (.A1(_10429_),
    .A2(_10571_),
    .ZN(_10573_));
 MUX2_X2 _19895_ (.A(_10572_),
    .B(_10573_),
    .S(_10444_),
    .Z(_10574_));
 AOI21_X4 _19896_ (.A(_10472_),
    .B1(_10448_),
    .B2(_10574_),
    .ZN(_10575_));
 NAND2_X4 _19897_ (.A1(_10558_),
    .A2(_10562_),
    .ZN(_10576_));
 AOI21_X2 _19898_ (.A(_10570_),
    .B1(_10575_),
    .B2(_10576_),
    .ZN(_10577_));
 BUF_X4 _19899_ (.A(_10494_),
    .Z(_10578_));
 AOI221_X2 _19900_ (.A(_10546_),
    .B1(_10563_),
    .B2(_10564_),
    .C1(_10577_),
    .C2(_10578_),
    .ZN(_10579_));
 NOR2_X2 _19901_ (.A1(_10568_),
    .A2(_10569_),
    .ZN(_10580_));
 BUF_X4 _19902_ (.A(_10580_),
    .Z(_10581_));
 BUF_X4 _19903_ (.A(_14862_),
    .Z(_10582_));
 BUF_X8 _19904_ (.A(_10558_),
    .Z(_10583_));
 BUF_X8 _19905_ (.A(_10562_),
    .Z(_10584_));
 NAND3_X4 _19906_ (.A1(_10471_),
    .A2(_10583_),
    .A3(_10584_),
    .ZN(_10585_));
 BUF_X8 _19907_ (.A(_10450_),
    .Z(_10586_));
 OAI221_X2 _19908_ (.A(_10500_),
    .B1(_10581_),
    .B2(_10582_),
    .C1(_10585_),
    .C2(_10586_),
    .ZN(_10587_));
 XNOR2_X2 _19909_ (.A(_06672_),
    .B(_10545_),
    .ZN(_10588_));
 BUF_X4 _19910_ (.A(_10588_),
    .Z(_10589_));
 NOR3_X4 _19911_ (.A1(_10494_),
    .A2(_10568_),
    .A3(_10569_),
    .ZN(_10590_));
 CLKBUF_X3 _19912_ (.A(_14868_),
    .Z(_10591_));
 INV_X2 _19913_ (.A(_10591_),
    .ZN(_10592_));
 AOI21_X2 _19914_ (.A(_10589_),
    .B1(_10590_),
    .B2(_10592_),
    .ZN(_10593_));
 AOI21_X2 _19915_ (.A(_10579_),
    .B1(_10587_),
    .B2(_10593_),
    .ZN(_10594_));
 BUF_X4 _19916_ (.A(_10533_),
    .Z(_10595_));
 BUF_X4 _19917_ (.A(_10546_),
    .Z(_10596_));
 BUF_X4 _19918_ (.A(_10596_),
    .Z(_10597_));
 BUF_X4 _19919_ (.A(_10597_),
    .Z(_10598_));
 BUF_X4 _19920_ (.A(_10576_),
    .Z(_10599_));
 CLKBUF_X3 _19921_ (.A(_10599_),
    .Z(_10600_));
 BUF_X4 _19922_ (.A(_14861_),
    .Z(_10601_));
 BUF_X16 _19923_ (.A(_10601_),
    .Z(_10602_));
 BUF_X4 _19924_ (.A(_10602_),
    .Z(_10603_));
 AOI22_X1 _19925_ (.A1(_14881_),
    .A2(_10600_),
    .B1(_10590_),
    .B2(_10603_),
    .ZN(_10604_));
 AOI21_X2 _19926_ (.A(_10595_),
    .B1(_10604_),
    .B2(_10598_),
    .ZN(_10605_));
 BUF_X4 _19927_ (.A(_10546_),
    .Z(_10606_));
 BUF_X4 _19928_ (.A(_10581_),
    .Z(_10607_));
 BUF_X2 split165 (.A(net985),
    .Z(net165));
 INV_X4 _19930_ (.A(net985),
    .ZN(_10609_));
 NOR2_X4 _19931_ (.A1(_10473_),
    .A2(_10496_),
    .ZN(_10610_));
 AOI22_X4 _19932_ (.A1(_10609_),
    .A2(_10497_),
    .B1(_10610_),
    .B2(_10452_),
    .ZN(_10611_));
 AOI21_X4 _19933_ (.A(_10606_),
    .B1(_10607_),
    .B2(_10611_),
    .ZN(_10612_));
 OAI21_X2 _19934_ (.A(_10494_),
    .B1(_10568_),
    .B2(_10569_),
    .ZN(_10613_));
 CLKBUF_X3 _19935_ (.A(_10613_),
    .Z(_10614_));
 BUF_X2 _19936_ (.A(_14860_),
    .Z(_10615_));
 CLKBUF_X3 _19937_ (.A(_10615_),
    .Z(_10616_));
 NAND2_X1 _19938_ (.A1(_10582_),
    .A2(_10607_),
    .ZN(_10617_));
 BUF_X8 _19939_ (.A(_10568_),
    .Z(_10618_));
 BUF_X8 _19940_ (.A(_10569_),
    .Z(_10619_));
 OAI21_X4 _19941_ (.A(_10473_),
    .B1(_10618_),
    .B2(_10619_),
    .ZN(_10620_));
 AND2_X1 _19942_ (.A1(_10617_),
    .A2(_10620_),
    .ZN(_10621_));
 BUF_X4 _19943_ (.A(_10578_),
    .Z(_10622_));
 BUF_X4 _19944_ (.A(_10622_),
    .Z(_10623_));
 OAI221_X2 _19945_ (.A(_10612_),
    .B1(_10614_),
    .B2(_10616_),
    .C1(_10621_),
    .C2(_10623_),
    .ZN(_10624_));
 AOI221_X2 _19946_ (.A(_10522_),
    .B1(_10534_),
    .B2(_10594_),
    .C1(_10605_),
    .C2(_10624_),
    .ZN(_10625_));
 XOR2_X2 _19947_ (.A(_06696_),
    .B(_10520_),
    .Z(_10626_));
 BUF_X4 _19948_ (.A(_10626_),
    .Z(_10627_));
 NAND2_X2 _19949_ (.A1(_10511_),
    .A2(_10627_),
    .ZN(_10628_));
 CLKBUF_X3 _19950_ (.A(_10588_),
    .Z(_10629_));
 NAND3_X1 _19951_ (.A1(_14858_),
    .A2(_10629_),
    .A3(_10600_),
    .ZN(_10630_));
 BUF_X4 _19952_ (.A(_10622_),
    .Z(_10631_));
 BUF_X4 _19953_ (.A(_10607_),
    .Z(_10632_));
 AOI21_X1 _19954_ (.A(_10631_),
    .B1(_10632_),
    .B2(_10609_),
    .ZN(_10633_));
 AOI21_X1 _19955_ (.A(_10595_),
    .B1(_10630_),
    .B2(_10633_),
    .ZN(_10634_));
 NOR2_X4 _19956_ (.A1(_10471_),
    .A2(_10495_),
    .ZN(_10635_));
 NAND2_X1 _19957_ (.A1(_10452_),
    .A2(_10635_),
    .ZN(_10636_));
 NAND2_X1 _19958_ (.A1(_10471_),
    .A2(_10496_),
    .ZN(_10637_));
 AND2_X1 _19959_ (.A1(_10576_),
    .A2(_10637_),
    .ZN(_10638_));
 AOI21_X4 _19960_ (.A(_10546_),
    .B1(_10636_),
    .B2(_10638_),
    .ZN(_10639_));
 INV_X2 _19961_ (.A(_14870_),
    .ZN(_10640_));
 NOR2_X2 _19962_ (.A1(_10640_),
    .A2(_10497_),
    .ZN(_10641_));
 NOR2_X4 _19963_ (.A1(_10495_),
    .A2(_10580_),
    .ZN(_10642_));
 AOI221_X2 _19964_ (.A(_10589_),
    .B1(_10607_),
    .B2(_10641_),
    .C1(_10642_),
    .C2(_10603_),
    .ZN(_10643_));
 OAI21_X1 _19965_ (.A(_10634_),
    .B1(_10639_),
    .B2(_10643_),
    .ZN(_10644_));
 XNOR2_X2 _19966_ (.A(_06687_),
    .B(_10531_),
    .ZN(_10645_));
 BUF_X4 _19967_ (.A(_10645_),
    .Z(_10646_));
 NOR2_X1 _19968_ (.A1(_10646_),
    .A2(_10589_),
    .ZN(_10647_));
 AOI21_X2 _19969_ (.A(net985),
    .B1(_10583_),
    .B2(_10584_),
    .ZN(_10648_));
 OAI21_X1 _19970_ (.A(_10623_),
    .B1(_10570_),
    .B2(_10648_),
    .ZN(_10649_));
 NAND3_X4 _19971_ (.A1(_10496_),
    .A2(_10583_),
    .A3(_10584_),
    .ZN(_10650_));
 INV_X1 _19972_ (.A(_10616_),
    .ZN(_10651_));
 OAI21_X1 _19973_ (.A(_10649_),
    .B1(_10650_),
    .B2(_10651_),
    .ZN(_10652_));
 NOR2_X2 _19974_ (.A1(_10645_),
    .A2(_10546_),
    .ZN(_10653_));
 BUF_X4 _19975_ (.A(_10581_),
    .Z(_10654_));
 BUF_X4 _19976_ (.A(_10654_),
    .Z(_10655_));
 NAND2_X4 _19977_ (.A1(_10473_),
    .A2(_10578_),
    .ZN(_10656_));
 BUF_X4 _19978_ (.A(_10497_),
    .Z(_10657_));
 NAND2_X1 _19979_ (.A1(_10592_),
    .A2(_10657_),
    .ZN(_10658_));
 AOI21_X1 _19980_ (.A(_10655_),
    .B1(_10656_),
    .B2(_10658_),
    .ZN(_10659_));
 BUF_X4 _19981_ (.A(_10576_),
    .Z(_10660_));
 AOI21_X2 _19982_ (.A(_10660_),
    .B1(_10578_),
    .B2(_10452_),
    .ZN(_10661_));
 NAND2_X1 _19983_ (.A1(_10603_),
    .A2(_10499_),
    .ZN(_10662_));
 AOI21_X1 _19984_ (.A(_10659_),
    .B1(_10661_),
    .B2(_10662_),
    .ZN(_10663_));
 AOI22_X1 _19985_ (.A1(_10647_),
    .A2(_10652_),
    .B1(_10653_),
    .B2(_10663_),
    .ZN(_10664_));
 AOI21_X1 _19986_ (.A(_10628_),
    .B1(_10644_),
    .B2(_10664_),
    .ZN(_10665_));
 NOR2_X4 _19987_ (.A1(_10511_),
    .A2(_10521_),
    .ZN(_10666_));
 INV_X1 _19988_ (.A(_10666_),
    .ZN(_10667_));
 BUF_X4 _19989_ (.A(_10452_),
    .Z(_10668_));
 NOR2_X1 _19990_ (.A1(_10668_),
    .A2(_10607_),
    .ZN(_10669_));
 OAI22_X1 _19991_ (.A1(net165),
    .A2(_10614_),
    .B1(_10637_),
    .B2(_10669_),
    .ZN(_10670_));
 NOR2_X1 _19992_ (.A1(_10582_),
    .A2(_10496_),
    .ZN(_10671_));
 AOI21_X4 _19993_ (.A(_10494_),
    .B1(_10448_),
    .B2(_10574_),
    .ZN(_10672_));
 NOR3_X2 _19994_ (.A1(_10576_),
    .A2(_10671_),
    .A3(_10672_),
    .ZN(_10673_));
 NOR2_X1 _19995_ (.A1(_10595_),
    .A2(_10673_),
    .ZN(_10674_));
 AOI22_X1 _19996_ (.A1(_10653_),
    .A2(_10670_),
    .B1(_10674_),
    .B2(_10639_),
    .ZN(_10675_));
 BUF_X2 split152 (.A(_15210_),
    .Z(net152));
 OAI21_X2 _19998_ (.A(_14874_),
    .B1(_10618_),
    .B2(_10619_),
    .ZN(_10677_));
 NAND2_X2 _19999_ (.A1(_10668_),
    .A2(_10654_),
    .ZN(_10678_));
 AND3_X1 _20000_ (.A1(_10631_),
    .A2(_10677_),
    .A3(_10678_),
    .ZN(_10679_));
 BUF_X4 _20001_ (.A(_10599_),
    .Z(_10680_));
 NOR2_X1 _20002_ (.A1(_14864_),
    .A2(_10680_),
    .ZN(_10681_));
 OAI21_X1 _20003_ (.A(_10646_),
    .B1(_10637_),
    .B2(_10681_),
    .ZN(_10682_));
 NOR3_X4 _20004_ (.A1(_10471_),
    .A2(_10618_),
    .A3(_10619_),
    .ZN(_10683_));
 OAI21_X1 _20005_ (.A(_10677_),
    .B1(_10599_),
    .B2(_10452_),
    .ZN(_10684_));
 AOI221_X1 _20006_ (.A(_10683_),
    .B1(_10684_),
    .B2(_10498_),
    .C1(_10602_),
    .C2(_10642_),
    .ZN(_10685_));
 BUF_X4 _20007_ (.A(_10646_),
    .Z(_10686_));
 OAI221_X1 _20008_ (.A(_10598_),
    .B1(_10679_),
    .B2(_10682_),
    .C1(_10685_),
    .C2(_10686_),
    .ZN(_10687_));
 AOI21_X1 _20009_ (.A(_10667_),
    .B1(_10675_),
    .B2(_10687_),
    .ZN(_10688_));
 CLKBUF_X3 _20010_ (.A(_10589_),
    .Z(_10689_));
 OAI21_X2 _20011_ (.A(_10473_),
    .B1(_10449_),
    .B2(_10445_),
    .ZN(_10690_));
 AND2_X1 _20012_ (.A1(_10581_),
    .A2(_10690_),
    .ZN(_10691_));
 OAI21_X1 _20013_ (.A(_10499_),
    .B1(_10655_),
    .B2(_10616_),
    .ZN(_10692_));
 NAND3_X2 _20014_ (.A1(_10602_),
    .A2(_10583_),
    .A3(_10584_),
    .ZN(_10693_));
 OAI21_X1 _20015_ (.A(_10693_),
    .B1(_10632_),
    .B2(_10591_),
    .ZN(_10694_));
 CLKBUF_X3 _20016_ (.A(_10657_),
    .Z(_10695_));
 OAI221_X1 _20017_ (.A(_10689_),
    .B1(_10691_),
    .B2(_10692_),
    .C1(_10694_),
    .C2(_10695_),
    .ZN(_10696_));
 NAND3_X4 _20018_ (.A1(_10574_),
    .A2(_10448_),
    .A3(_10471_),
    .ZN(_10697_));
 NAND2_X1 _20019_ (.A1(_10656_),
    .A2(_10697_),
    .ZN(_10698_));
 XNOR2_X1 _20020_ (.A(_10632_),
    .B(_10698_),
    .ZN(_10699_));
 OAI21_X1 _20021_ (.A(_10696_),
    .B1(_10699_),
    .B2(_10689_),
    .ZN(_10700_));
 NOR2_X4 _20022_ (.A1(_10511_),
    .A2(_10626_),
    .ZN(_10701_));
 NAND2_X1 _20023_ (.A1(_10534_),
    .A2(_10701_),
    .ZN(_10702_));
 NAND2_X2 _20024_ (.A1(_10521_),
    .A2(_10546_),
    .ZN(_10703_));
 NOR2_X2 _20025_ (.A1(_10602_),
    .A2(_10578_),
    .ZN(_10704_));
 NAND2_X2 _20026_ (.A1(net988),
    .A2(_10581_),
    .ZN(_10705_));
 NAND2_X1 _20027_ (.A1(net987),
    .A2(_10497_),
    .ZN(_10706_));
 INV_X4 _20028_ (.A(_10601_),
    .ZN(_10707_));
 NOR3_X4 _20029_ (.A1(_10707_),
    .A2(_10618_),
    .A3(_10619_),
    .ZN(_10708_));
 AOI221_X1 _20030_ (.A(_10703_),
    .B1(_10704_),
    .B2(_10705_),
    .C1(_10706_),
    .C2(_10708_),
    .ZN(_10709_));
 NAND2_X1 _20031_ (.A1(_10591_),
    .A2(_10590_),
    .ZN(_10710_));
 NOR3_X4 _20032_ (.A1(_10495_),
    .A2(_10568_),
    .A3(_10569_),
    .ZN(_10711_));
 NOR2_X2 _20033_ (.A1(_10563_),
    .A2(_10711_),
    .ZN(_10712_));
 OAI221_X1 _20034_ (.A(_10710_),
    .B1(_10712_),
    .B2(_10651_),
    .C1(_10614_),
    .C2(_10603_),
    .ZN(_10713_));
 NOR2_X2 _20035_ (.A1(_10627_),
    .A2(_10606_),
    .ZN(_10714_));
 AOI21_X1 _20036_ (.A(_10709_),
    .B1(_10713_),
    .B2(_10714_),
    .ZN(_10715_));
 XNOR2_X2 _20037_ (.A(_06710_),
    .B(_10510_),
    .ZN(_10716_));
 NAND2_X1 _20038_ (.A1(_10716_),
    .A2(_10646_),
    .ZN(_10717_));
 OAI22_X1 _20039_ (.A1(_10700_),
    .A2(_10702_),
    .B1(_10715_),
    .B2(_10717_),
    .ZN(_10718_));
 NOR4_X1 _20040_ (.A1(_10718_),
    .A2(_10665_),
    .A3(_10688_),
    .A4(_10625_),
    .ZN(_00048_));
 CLKBUF_X3 _20041_ (.A(_10686_),
    .Z(_10719_));
 NAND2_X2 _20042_ (.A1(_10626_),
    .A2(_10588_),
    .ZN(_10720_));
 AND2_X1 _20043_ (.A1(_10660_),
    .A2(_10690_),
    .ZN(_10721_));
 NOR2_X1 _20044_ (.A1(_14876_),
    .A2(_10721_),
    .ZN(_10722_));
 AOI21_X4 _20045_ (.A(_10602_),
    .B1(_10583_),
    .B2(_10584_),
    .ZN(_10723_));
 NOR2_X1 _20046_ (.A1(_10609_),
    .A2(_10660_),
    .ZN(_10724_));
 NOR3_X1 _20047_ (.A1(_14883_),
    .A2(_10723_),
    .A3(_10724_),
    .ZN(_10725_));
 NOR3_X1 _20048_ (.A1(_10720_),
    .A2(_10722_),
    .A3(_10725_),
    .ZN(_10726_));
 NAND3_X4 _20049_ (.A1(_10473_),
    .A2(_10583_),
    .A3(_10584_),
    .ZN(_10727_));
 NOR2_X2 _20050_ (.A1(_10586_),
    .A2(_10727_),
    .ZN(_10728_));
 NAND2_X2 _20051_ (.A1(_10626_),
    .A2(_10546_),
    .ZN(_10729_));
 INV_X2 _20052_ (.A(_14874_),
    .ZN(_10730_));
 AOI21_X1 _20053_ (.A(_10730_),
    .B1(_10583_),
    .B2(_10584_),
    .ZN(_10731_));
 OAI22_X1 _20054_ (.A1(_14864_),
    .A2(_10614_),
    .B1(_10731_),
    .B2(_10623_),
    .ZN(_10732_));
 NOR3_X2 _20055_ (.A1(_10728_),
    .A2(_10729_),
    .A3(_10732_),
    .ZN(_10733_));
 NAND2_X1 _20056_ (.A1(_10597_),
    .A2(_10563_),
    .ZN(_10734_));
 BUF_X16 _20057_ (.A(_10586_),
    .Z(_10735_));
 NAND3_X1 _20058_ (.A1(_10735_),
    .A2(_10629_),
    .A3(_10655_),
    .ZN(_10736_));
 AOI21_X1 _20059_ (.A(_14867_),
    .B1(_10734_),
    .B2(_10736_),
    .ZN(_10737_));
 NAND3_X1 _20060_ (.A1(_10609_),
    .A2(_10596_),
    .A3(_10654_),
    .ZN(_10738_));
 OAI21_X1 _20061_ (.A(_10680_),
    .B1(_10589_),
    .B2(_10707_),
    .ZN(_10739_));
 AOI21_X1 _20062_ (.A(_10499_),
    .B1(_10738_),
    .B2(_10739_),
    .ZN(_10740_));
 BUF_X16 _20063_ (.A(_10735_),
    .Z(_14859_));
 AOI22_X1 _20064_ (.A1(_10501_),
    .A2(_10589_),
    .B1(_10563_),
    .B2(_14858_),
    .ZN(_10741_));
 NAND2_X1 _20065_ (.A1(_10606_),
    .A2(_10655_),
    .ZN(_10742_));
 NAND2_X2 _20066_ (.A1(_10473_),
    .A2(_10496_),
    .ZN(_10743_));
 OAI22_X1 _20067_ (.A1(_14859_),
    .A2(_10741_),
    .B1(_10742_),
    .B2(_10743_),
    .ZN(_10744_));
 NOR4_X2 _20068_ (.A1(_10627_),
    .A2(_10737_),
    .A3(_10740_),
    .A4(_10744_),
    .ZN(_10745_));
 NOR4_X2 _20069_ (.A1(_10719_),
    .A2(_10726_),
    .A3(_10733_),
    .A4(_10745_),
    .ZN(_10746_));
 NOR2_X1 _20070_ (.A1(_10707_),
    .A2(_10622_),
    .ZN(_10747_));
 NOR2_X1 _20071_ (.A1(_10730_),
    .A2(_10657_),
    .ZN(_10748_));
 OAI21_X1 _20072_ (.A(_10680_),
    .B1(_10747_),
    .B2(_10748_),
    .ZN(_10749_));
 OAI22_X2 _20073_ (.A1(net165),
    .A2(_10650_),
    .B1(_10712_),
    .B2(_10735_),
    .ZN(_10750_));
 AOI221_X2 _20074_ (.A(_10522_),
    .B1(_10612_),
    .B2(_10749_),
    .C1(_10750_),
    .C2(_10598_),
    .ZN(_10751_));
 OAI222_X2 _20075_ (.A1(_14864_),
    .A2(_10620_),
    .B1(_10712_),
    .B2(_14867_),
    .C1(_10650_),
    .C2(_10707_),
    .ZN(_10752_));
 NOR3_X1 _20076_ (.A1(_10598_),
    .A2(_10628_),
    .A3(_10752_),
    .ZN(_10753_));
 NOR3_X2 _20077_ (.A1(_10473_),
    .A2(_10618_),
    .A3(_10619_),
    .ZN(_10754_));
 NOR3_X1 _20078_ (.A1(_10631_),
    .A2(_10754_),
    .A3(_10648_),
    .ZN(_10755_));
 OAI21_X4 _20079_ (.A(_10707_),
    .B1(_10618_),
    .B2(_10619_),
    .ZN(_10756_));
 OAI21_X1 _20080_ (.A(_10756_),
    .B1(_10600_),
    .B2(_10616_),
    .ZN(_10757_));
 AOI21_X1 _20081_ (.A(_10755_),
    .B1(_10757_),
    .B2(_14876_),
    .ZN(_10758_));
 NAND3_X1 _20082_ (.A1(_10511_),
    .A2(_10627_),
    .A3(_10598_),
    .ZN(_10759_));
 OAI22_X1 _20083_ (.A1(_10716_),
    .A2(_10719_),
    .B1(_10758_),
    .B2(_10759_),
    .ZN(_10760_));
 NOR3_X2 _20084_ (.A1(_10751_),
    .A2(_10753_),
    .A3(_10760_),
    .ZN(_10761_));
 OAI221_X2 _20085_ (.A(_10654_),
    .B1(_10656_),
    .B2(_10586_),
    .C1(_10500_),
    .C2(_10592_),
    .ZN(_10762_));
 INV_X1 _20086_ (.A(_14884_),
    .ZN(_10763_));
 BUF_X4 _20087_ (.A(_10680_),
    .Z(_10764_));
 NAND3_X1 _20088_ (.A1(_10763_),
    .A2(_10719_),
    .A3(_10764_),
    .ZN(_10765_));
 NAND3_X1 _20089_ (.A1(_10714_),
    .A2(_10762_),
    .A3(_10765_),
    .ZN(_10766_));
 INV_X1 _20090_ (.A(_10703_),
    .ZN(_10767_));
 OAI21_X1 _20091_ (.A(_10631_),
    .B1(_10648_),
    .B2(_10683_),
    .ZN(_10768_));
 XNOR2_X2 _20092_ (.A(net987),
    .B(_10654_),
    .ZN(_10769_));
 OAI211_X2 _20093_ (.A(_10686_),
    .B(_10768_),
    .C1(_10769_),
    .C2(_14876_),
    .ZN(_10770_));
 NAND2_X1 _20094_ (.A1(_14864_),
    .A2(_10764_),
    .ZN(_10771_));
 XNOR2_X1 _20095_ (.A(_14867_),
    .B(_10498_),
    .ZN(_10772_));
 AOI21_X1 _20096_ (.A(_10610_),
    .B1(_14883_),
    .B2(_10616_),
    .ZN(_10773_));
 OAI221_X1 _20097_ (.A(_10534_),
    .B1(_10771_),
    .B2(_10772_),
    .C1(_10773_),
    .C2(_10764_),
    .ZN(_10774_));
 NAND3_X1 _20098_ (.A1(_10767_),
    .A2(_10770_),
    .A3(_10774_),
    .ZN(_10775_));
 NAND3_X1 _20099_ (.A1(_10716_),
    .A2(_10766_),
    .A3(_10775_),
    .ZN(_10776_));
 OAI21_X1 _20100_ (.A(_10756_),
    .B1(_10727_),
    .B2(_10735_),
    .ZN(_10777_));
 AOI221_X2 _20101_ (.A(_10533_),
    .B1(_10590_),
    .B2(_14858_),
    .C1(_10777_),
    .C2(_10631_),
    .ZN(_10778_));
 INV_X1 _20102_ (.A(_10768_),
    .ZN(_10779_));
 NOR2_X1 _20103_ (.A1(_10616_),
    .A2(_10680_),
    .ZN(_10780_));
 NOR2_X2 _20104_ (.A1(net989),
    .A2(_10581_),
    .ZN(_10781_));
 NOR3_X1 _20105_ (.A1(_10623_),
    .A2(_10780_),
    .A3(_10781_),
    .ZN(_10782_));
 NOR3_X1 _20106_ (.A1(_10719_),
    .A2(_10779_),
    .A3(_10782_),
    .ZN(_10783_));
 NAND3_X1 _20107_ (.A1(_10695_),
    .A2(_10585_),
    .A3(_10756_),
    .ZN(_10784_));
 AOI21_X1 _20108_ (.A(_10570_),
    .B1(_10600_),
    .B2(_10616_),
    .ZN(_10785_));
 NAND2_X1 _20109_ (.A1(_14876_),
    .A2(_10785_),
    .ZN(_10786_));
 AOI21_X1 _20110_ (.A(_10686_),
    .B1(_10784_),
    .B2(_10786_),
    .ZN(_10787_));
 CLKBUF_X3 _20111_ (.A(_10660_),
    .Z(_10788_));
 NAND2_X1 _20112_ (.A1(_10788_),
    .A2(_10690_),
    .ZN(_10789_));
 AOI21_X1 _20113_ (.A(_10500_),
    .B1(_10654_),
    .B2(_10582_),
    .ZN(_10790_));
 AOI21_X2 _20114_ (.A(_10723_),
    .B1(_10607_),
    .B2(net166),
    .ZN(_10791_));
 AOI221_X2 _20115_ (.A(_10533_),
    .B1(_10789_),
    .B2(_10790_),
    .C1(_10791_),
    .C2(_10501_),
    .ZN(_10792_));
 OAI33_X1 _20116_ (.A1(_10720_),
    .A2(_10778_),
    .A3(_10783_),
    .B1(_10792_),
    .B2(_10787_),
    .B3(_10729_),
    .ZN(_10793_));
 OAI22_X2 _20117_ (.A1(_10746_),
    .A2(_10761_),
    .B1(_10793_),
    .B2(_10776_),
    .ZN(_00049_));
 AND2_X1 _20118_ (.A1(_10662_),
    .A2(_10661_),
    .ZN(_10794_));
 OAI21_X1 _20119_ (.A(_10629_),
    .B1(_10632_),
    .B2(_10611_),
    .ZN(_10795_));
 NOR3_X1 _20120_ (.A1(_10627_),
    .A2(_10794_),
    .A3(_10795_),
    .ZN(_10796_));
 NOR3_X4 _20121_ (.A1(net848),
    .A2(_10568_),
    .A3(_10569_),
    .ZN(_10797_));
 NOR3_X1 _20122_ (.A1(_10501_),
    .A2(_10648_),
    .A3(_10797_),
    .ZN(_10798_));
 MUX2_X1 _20123_ (.A(_10564_),
    .B(_14867_),
    .S(_10599_),
    .Z(_10799_));
 AOI21_X1 _20124_ (.A(_10798_),
    .B1(_10799_),
    .B2(_10623_),
    .ZN(_10800_));
 NOR2_X1 _20125_ (.A1(_10729_),
    .A2(_10800_),
    .ZN(_10801_));
 MUX2_X1 _20126_ (.A(_14874_),
    .B(_14865_),
    .S(_10494_),
    .Z(_10802_));
 INV_X1 _20127_ (.A(_10802_),
    .ZN(_10803_));
 AOI221_X1 _20128_ (.A(_10703_),
    .B1(_10743_),
    .B2(_10781_),
    .C1(_10803_),
    .C2(_10581_),
    .ZN(_10804_));
 AOI21_X1 _20129_ (.A(_10496_),
    .B1(_10576_),
    .B2(_10451_),
    .ZN(_10805_));
 NAND3_X2 _20130_ (.A1(_10564_),
    .A2(_10558_),
    .A3(_10562_),
    .ZN(_10806_));
 AOI221_X1 _20131_ (.A(_10720_),
    .B1(_10805_),
    .B2(_10806_),
    .C1(_10497_),
    .C2(_10609_),
    .ZN(_10807_));
 OR3_X1 _20132_ (.A1(_10717_),
    .A2(_10804_),
    .A3(_10807_),
    .ZN(_10808_));
 OR3_X1 _20133_ (.A1(_10796_),
    .A2(_10801_),
    .A3(_10808_),
    .ZN(_10809_));
 INV_X1 _20134_ (.A(_14888_),
    .ZN(_10810_));
 AOI221_X1 _20135_ (.A(_10703_),
    .B1(_10743_),
    .B2(_10781_),
    .C1(_10655_),
    .C2(_10810_),
    .ZN(_10811_));
 NOR3_X1 _20136_ (.A1(_10716_),
    .A2(_10534_),
    .A3(_10811_),
    .ZN(_10812_));
 CLKBUF_X3 _20137_ (.A(_10655_),
    .Z(_10813_));
 NOR2_X1 _20138_ (.A1(_14879_),
    .A2(_10813_),
    .ZN(_10814_));
 NAND2_X1 _20139_ (.A1(_10497_),
    .A2(_10575_),
    .ZN(_10815_));
 AOI21_X1 _20140_ (.A(_10814_),
    .B1(_10815_),
    .B2(_10813_),
    .ZN(_10816_));
 NAND2_X1 _20141_ (.A1(_10521_),
    .A2(_10588_),
    .ZN(_10817_));
 AOI21_X1 _20142_ (.A(_10597_),
    .B1(_10813_),
    .B2(_10763_),
    .ZN(_10818_));
 OAI21_X1 _20143_ (.A(_10697_),
    .B1(_10695_),
    .B2(_14859_),
    .ZN(_10819_));
 OAI21_X1 _20144_ (.A(_10818_),
    .B1(_10819_),
    .B2(_10813_),
    .ZN(_10820_));
 NAND3_X4 _20145_ (.A1(_10615_),
    .A2(_10583_),
    .A3(_10584_),
    .ZN(_10821_));
 NAND3_X1 _20146_ (.A1(_10695_),
    .A2(_10756_),
    .A3(_10821_),
    .ZN(_10822_));
 MUX2_X1 _20147_ (.A(_10591_),
    .B(_10735_),
    .S(_10655_),
    .Z(_10823_));
 OAI21_X1 _20148_ (.A(_10822_),
    .B1(_10823_),
    .B2(_14883_),
    .ZN(_10824_));
 OAI21_X1 _20149_ (.A(_10820_),
    .B1(_10824_),
    .B2(_10689_),
    .ZN(_10825_));
 OAI221_X1 _20150_ (.A(_10812_),
    .B1(_10816_),
    .B2(_10817_),
    .C1(_10825_),
    .C2(_10521_),
    .ZN(_10826_));
 NAND2_X1 _20151_ (.A1(_10620_),
    .A2(_10585_),
    .ZN(_10827_));
 AOI221_X1 _20152_ (.A(_10817_),
    .B1(_10827_),
    .B2(_10672_),
    .C1(_10642_),
    .C2(_10730_),
    .ZN(_10828_));
 NOR3_X1 _20153_ (.A1(_10511_),
    .A2(_10719_),
    .A3(_10828_),
    .ZN(_10829_));
 OAI21_X2 _20154_ (.A(_10640_),
    .B1(_10568_),
    .B2(_10569_),
    .ZN(_10830_));
 AND2_X1 _20155_ (.A1(_10585_),
    .A2(_10830_),
    .ZN(_10831_));
 AOI21_X1 _20156_ (.A(_10797_),
    .B1(_10680_),
    .B2(_10668_),
    .ZN(_10832_));
 MUX2_X1 _20157_ (.A(_10831_),
    .B(_10832_),
    .S(_10499_),
    .Z(_10833_));
 OAI21_X1 _20158_ (.A(_10817_),
    .B1(_10729_),
    .B2(_10833_),
    .ZN(_10834_));
 AND2_X1 _20159_ (.A1(_10620_),
    .A2(_10693_),
    .ZN(_10835_));
 NOR2_X1 _20160_ (.A1(_14883_),
    .A2(_10835_),
    .ZN(_10836_));
 NAND2_X1 _20161_ (.A1(_10582_),
    .A2(_10599_),
    .ZN(_10837_));
 AOI21_X1 _20162_ (.A(_10623_),
    .B1(_10837_),
    .B2(_10705_),
    .ZN(_10838_));
 NOR3_X1 _20163_ (.A1(_10695_),
    .A2(_10754_),
    .A3(_10723_),
    .ZN(_10839_));
 AOI21_X1 _20164_ (.A(_10631_),
    .B1(_10806_),
    .B2(_10756_),
    .ZN(_10840_));
 OAI33_X1 _20165_ (.A1(_10627_),
    .A2(_10836_),
    .A3(_10838_),
    .B1(_10839_),
    .B2(_10840_),
    .B3(_10597_),
    .ZN(_10841_));
 OAI21_X1 _20166_ (.A(_10829_),
    .B1(_10834_),
    .B2(_10841_),
    .ZN(_10842_));
 NOR2_X1 _20167_ (.A1(_10716_),
    .A2(_10719_),
    .ZN(_10843_));
 OR2_X1 _20168_ (.A1(_10654_),
    .A2(_10690_),
    .ZN(_10844_));
 NAND3_X2 _20169_ (.A1(_10591_),
    .A2(_10583_),
    .A3(_10584_),
    .ZN(_10845_));
 AND2_X1 _20170_ (.A1(_10497_),
    .A2(_10845_),
    .ZN(_10846_));
 NOR2_X2 _20171_ (.A1(_10582_),
    .A2(net985),
    .ZN(_10847_));
 AOI21_X1 _20172_ (.A(_10728_),
    .B1(_10847_),
    .B2(_10788_),
    .ZN(_10848_));
 AOI221_X2 _20173_ (.A(_10589_),
    .B1(_10844_),
    .B2(_10846_),
    .C1(_10848_),
    .C2(_10631_),
    .ZN(_10849_));
 NAND3_X1 _20174_ (.A1(_10501_),
    .A2(_10756_),
    .A3(_10821_),
    .ZN(_10850_));
 OAI21_X4 _20175_ (.A(_10496_),
    .B1(_10618_),
    .B2(_10619_),
    .ZN(_10851_));
 OAI21_X1 _20176_ (.A(_10850_),
    .B1(_10851_),
    .B2(_10609_),
    .ZN(_10852_));
 OAI21_X1 _20177_ (.A(_10521_),
    .B1(_10598_),
    .B2(_10852_),
    .ZN(_10853_));
 NAND3_X1 _20178_ (.A1(_10668_),
    .A2(_10501_),
    .A3(_10620_),
    .ZN(_10854_));
 NAND2_X1 _20179_ (.A1(_10735_),
    .A2(_10788_),
    .ZN(_10855_));
 MUX2_X1 _20180_ (.A(_10500_),
    .B(_10599_),
    .S(_10452_),
    .Z(_10856_));
 OAI221_X1 _20181_ (.A(_10854_),
    .B1(_10855_),
    .B2(_10635_),
    .C1(_10707_),
    .C2(_10856_),
    .ZN(_10857_));
 NAND2_X1 _20182_ (.A1(_10500_),
    .A2(_10575_),
    .ZN(_10858_));
 NOR2_X1 _20183_ (.A1(_10655_),
    .A2(_10704_),
    .ZN(_10859_));
 AOI22_X1 _20184_ (.A1(_14881_),
    .A2(_10632_),
    .B1(_10858_),
    .B2(_10859_),
    .ZN(_10860_));
 MUX2_X1 _20185_ (.A(_10857_),
    .B(_10860_),
    .S(_10689_),
    .Z(_10861_));
 OAI221_X1 _20186_ (.A(_10843_),
    .B1(_10849_),
    .B2(_10853_),
    .C1(_10861_),
    .C2(_10521_),
    .ZN(_10862_));
 AND4_X1 _20187_ (.A1(_10809_),
    .A2(_10826_),
    .A3(_10842_),
    .A4(_10862_),
    .ZN(_00050_));
 OR2_X1 _20188_ (.A1(_14862_),
    .A2(_14865_),
    .ZN(_10863_));
 MUX2_X1 _20189_ (.A(_10564_),
    .B(_10863_),
    .S(_10494_),
    .Z(_10864_));
 AOI211_X2 _20190_ (.A(_10532_),
    .B(_10546_),
    .C1(_10660_),
    .C2(_10864_),
    .ZN(_10865_));
 AOI21_X1 _20191_ (.A(_10521_),
    .B1(_10762_),
    .B2(_10865_),
    .ZN(_10866_));
 AOI21_X1 _20192_ (.A(_14858_),
    .B1(_10622_),
    .B2(_10705_),
    .ZN(_10867_));
 OAI221_X1 _20193_ (.A(_10653_),
    .B1(_10650_),
    .B2(net987),
    .C1(_10616_),
    .C2(_10613_),
    .ZN(_10868_));
 OAI21_X1 _20194_ (.A(_10622_),
    .B1(_10532_),
    .B2(_10585_),
    .ZN(_10869_));
 OAI21_X1 _20195_ (.A(_10830_),
    .B1(_10576_),
    .B2(_10601_),
    .ZN(_10870_));
 AOI21_X1 _20196_ (.A(_10869_),
    .B1(_10870_),
    .B2(_10533_),
    .ZN(_10871_));
 OAI22_X1 _20197_ (.A1(net166),
    .A2(_10599_),
    .B1(_10620_),
    .B2(_10645_),
    .ZN(_10872_));
 OAI21_X1 _20198_ (.A(_10606_),
    .B1(_10872_),
    .B2(_10501_),
    .ZN(_10873_));
 OAI221_X1 _20199_ (.A(_10866_),
    .B1(_10867_),
    .B2(_10868_),
    .C1(_10871_),
    .C2(_10873_),
    .ZN(_10874_));
 NAND3_X4 _20200_ (.A1(_10494_),
    .A2(_10558_),
    .A3(_10562_),
    .ZN(_10875_));
 NAND2_X1 _20201_ (.A1(_10851_),
    .A2(_10875_),
    .ZN(_10876_));
 NOR2_X1 _20202_ (.A1(_10640_),
    .A2(_10876_),
    .ZN(_10877_));
 OAI21_X1 _20203_ (.A(_10533_),
    .B1(_10788_),
    .B2(_10656_),
    .ZN(_10878_));
 OAI21_X1 _20204_ (.A(_10498_),
    .B1(_10731_),
    .B2(_10683_),
    .ZN(_10879_));
 OAI21_X1 _20205_ (.A(_10847_),
    .B1(_10619_),
    .B2(_10618_),
    .ZN(_10880_));
 OAI21_X1 _20206_ (.A(_10880_),
    .B1(_10599_),
    .B2(_10602_),
    .ZN(_10881_));
 OAI21_X1 _20207_ (.A(_10879_),
    .B1(_10881_),
    .B2(_10499_),
    .ZN(_10882_));
 OAI221_X1 _20208_ (.A(_10714_),
    .B1(_10877_),
    .B2(_10878_),
    .C1(_10882_),
    .C2(_10595_),
    .ZN(_10883_));
 NAND2_X1 _20209_ (.A1(_10735_),
    .A2(_10711_),
    .ZN(_10884_));
 NOR3_X1 _20210_ (.A1(_10591_),
    .A2(_10618_),
    .A3(_10619_),
    .ZN(_10885_));
 OAI21_X1 _20211_ (.A(_10657_),
    .B1(_10723_),
    .B2(_10885_),
    .ZN(_10886_));
 AOI21_X1 _20212_ (.A(_10533_),
    .B1(_10884_),
    .B2(_10886_),
    .ZN(_10887_));
 NAND3_X1 _20213_ (.A1(_10707_),
    .A2(_10533_),
    .A3(_10654_),
    .ZN(_10888_));
 AOI21_X1 _20214_ (.A(_10657_),
    .B1(_10837_),
    .B2(_10888_),
    .ZN(_10889_));
 OAI21_X1 _20215_ (.A(_10767_),
    .B1(_10887_),
    .B2(_10889_),
    .ZN(_10890_));
 AND4_X1 _20216_ (.A1(_10716_),
    .A2(_10874_),
    .A3(_10883_),
    .A4(_10890_),
    .ZN(_10891_));
 NOR2_X2 _20217_ (.A1(_10532_),
    .A2(_10596_),
    .ZN(_10892_));
 AND4_X1 _20218_ (.A1(_10614_),
    .A2(_10697_),
    .A3(_10743_),
    .A4(_10892_),
    .ZN(_10893_));
 NOR2_X2 _20219_ (.A1(_10532_),
    .A2(_10588_),
    .ZN(_10894_));
 AOI21_X1 _20220_ (.A(_10501_),
    .B1(_10806_),
    .B2(_10677_),
    .ZN(_10895_));
 AOI21_X2 _20221_ (.A(_10708_),
    .B1(_10788_),
    .B2(_10735_),
    .ZN(_10896_));
 AOI21_X1 _20222_ (.A(_10895_),
    .B1(_10896_),
    .B2(_10623_),
    .ZN(_10897_));
 AOI21_X1 _20223_ (.A(_10893_),
    .B1(_10894_),
    .B2(_10897_),
    .ZN(_10898_));
 OAI221_X1 _20224_ (.A(_10710_),
    .B1(_10835_),
    .B2(_10657_),
    .C1(_10655_),
    .C2(_10697_),
    .ZN(_10899_));
 OAI221_X1 _20225_ (.A(_10629_),
    .B1(_10614_),
    .B2(_10592_),
    .C1(_10650_),
    .C2(_10603_),
    .ZN(_10900_));
 AOI22_X1 _20226_ (.A1(_14858_),
    .A2(_10563_),
    .B1(_10635_),
    .B2(_10607_),
    .ZN(_10901_));
 NOR2_X1 _20227_ (.A1(_14859_),
    .A2(_10901_),
    .ZN(_10902_));
 OAI221_X1 _20228_ (.A(_10595_),
    .B1(_10629_),
    .B2(_10899_),
    .C1(_10900_),
    .C2(_10902_),
    .ZN(_10903_));
 AOI21_X1 _20229_ (.A(_10628_),
    .B1(_10898_),
    .B2(_10903_),
    .ZN(_10904_));
 AOI21_X1 _20230_ (.A(_10708_),
    .B1(_10600_),
    .B2(_10730_),
    .ZN(_10905_));
 NAND2_X1 _20231_ (.A1(_14876_),
    .A2(_10905_),
    .ZN(_10906_));
 NAND2_X1 _20232_ (.A1(_10609_),
    .A2(_10788_),
    .ZN(_10907_));
 NAND3_X1 _20233_ (.A1(_10695_),
    .A2(_10907_),
    .A3(_10705_),
    .ZN(_10908_));
 AOI21_X1 _20234_ (.A(_10686_),
    .B1(_10906_),
    .B2(_10908_),
    .ZN(_10909_));
 NAND2_X1 _20235_ (.A1(_10616_),
    .A2(_10600_),
    .ZN(_10910_));
 NAND3_X1 _20236_ (.A1(_14876_),
    .A2(_10845_),
    .A3(_10910_),
    .ZN(_10911_));
 OAI21_X1 _20237_ (.A(_10695_),
    .B1(_10683_),
    .B2(_10723_),
    .ZN(_10912_));
 AOI21_X1 _20238_ (.A(_10686_),
    .B1(_10911_),
    .B2(_10912_),
    .ZN(_10913_));
 OAI21_X1 _20239_ (.A(_10598_),
    .B1(_10656_),
    .B2(_10534_),
    .ZN(_10914_));
 OAI22_X2 _20240_ (.A1(_10598_),
    .A2(_10909_),
    .B1(_10913_),
    .B2(_10914_),
    .ZN(_10915_));
 NAND2_X1 _20241_ (.A1(_10668_),
    .A2(_10589_),
    .ZN(_10916_));
 NOR2_X1 _20242_ (.A1(_10602_),
    .A2(_10498_),
    .ZN(_10917_));
 NOR2_X1 _20243_ (.A1(_10754_),
    .A2(_10917_),
    .ZN(_10918_));
 AOI22_X1 _20244_ (.A1(_10735_),
    .A2(_10606_),
    .B1(_10697_),
    .B2(_10622_),
    .ZN(_10919_));
 OAI221_X1 _20245_ (.A(_10686_),
    .B1(_10916_),
    .B2(_10918_),
    .C1(_10919_),
    .C2(_10600_),
    .ZN(_10920_));
 MUX2_X1 _20246_ (.A(_10668_),
    .B(_10622_),
    .S(_10596_),
    .Z(_10921_));
 OAI22_X1 _20247_ (.A1(_10597_),
    .A2(_10706_),
    .B1(_10921_),
    .B2(_10603_),
    .ZN(_10922_));
 AOI21_X1 _20248_ (.A(_10920_),
    .B1(_10922_),
    .B2(_10764_),
    .ZN(_10923_));
 NOR2_X1 _20249_ (.A1(_10522_),
    .A2(_10923_),
    .ZN(_10924_));
 AOI211_X2 _20250_ (.A(_10891_),
    .B(_10904_),
    .C1(_10915_),
    .C2(_10924_),
    .ZN(_00051_));
 NAND2_X1 _20251_ (.A1(_10668_),
    .A2(_10754_),
    .ZN(_10925_));
 NAND3_X1 _20252_ (.A1(_10646_),
    .A2(_10788_),
    .A3(_10635_),
    .ZN(_10926_));
 NAND4_X1 _20253_ (.A1(_10597_),
    .A2(_10925_),
    .A3(_10701_),
    .A4(_10926_),
    .ZN(_10927_));
 OAI21_X1 _20254_ (.A(_10650_),
    .B1(_10614_),
    .B2(_10646_),
    .ZN(_10928_));
 OAI21_X1 _20255_ (.A(_10830_),
    .B1(_10764_),
    .B2(_10646_),
    .ZN(_10929_));
 AOI221_X1 _20256_ (.A(_10927_),
    .B1(_10928_),
    .B2(_14859_),
    .C1(_14883_),
    .C2(_10929_),
    .ZN(_10930_));
 MUX2_X1 _20257_ (.A(_10582_),
    .B(_10690_),
    .S(_10660_),
    .Z(_10931_));
 NAND3_X1 _20258_ (.A1(_10498_),
    .A2(_10533_),
    .A3(_10596_),
    .ZN(_10932_));
 AOI22_X1 _20259_ (.A1(_10730_),
    .A2(_10590_),
    .B1(_10585_),
    .B2(_10622_),
    .ZN(_10933_));
 NAND2_X2 _20260_ (.A1(_10645_),
    .A2(_10588_),
    .ZN(_10934_));
 OAI221_X2 _20261_ (.A(_10666_),
    .B1(_10931_),
    .B2(_10932_),
    .C1(_10933_),
    .C2(_10934_),
    .ZN(_10935_));
 NAND2_X2 _20262_ (.A1(_10645_),
    .A2(_10546_),
    .ZN(_10936_));
 AOI21_X1 _20263_ (.A(_10936_),
    .B1(_10769_),
    .B2(_10499_),
    .ZN(_10937_));
 NAND3_X1 _20264_ (.A1(_10501_),
    .A2(_10907_),
    .A3(_10821_),
    .ZN(_10938_));
 MUX2_X1 _20265_ (.A(_10707_),
    .B(net165),
    .S(_10500_),
    .Z(_10939_));
 AOI21_X1 _20266_ (.A(_10646_),
    .B1(_10632_),
    .B2(_10939_),
    .ZN(_10940_));
 AOI221_X2 _20267_ (.A(_10935_),
    .B1(_10937_),
    .B2(_10938_),
    .C1(_10639_),
    .C2(_10940_),
    .ZN(_10941_));
 NOR2_X1 _20268_ (.A1(_10930_),
    .A2(_10941_),
    .ZN(_10942_));
 NAND3_X1 _20269_ (.A1(_10680_),
    .A2(_10858_),
    .A3(_10706_),
    .ZN(_10943_));
 AOI21_X1 _20270_ (.A(_10589_),
    .B1(_10607_),
    .B2(net986),
    .ZN(_10944_));
 NOR2_X1 _20271_ (.A1(_10616_),
    .A2(_10498_),
    .ZN(_10945_));
 OAI21_X1 _20272_ (.A(_10680_),
    .B1(_10672_),
    .B2(_10945_),
    .ZN(_10946_));
 AOI221_X2 _20273_ (.A(_10595_),
    .B1(_10944_),
    .B2(_10943_),
    .C1(_10946_),
    .C2(_10612_),
    .ZN(_10947_));
 NAND2_X2 _20274_ (.A1(_10576_),
    .A2(_10575_),
    .ZN(_10948_));
 NOR2_X1 _20275_ (.A1(_10596_),
    .A2(_10797_),
    .ZN(_10949_));
 NAND2_X1 _20276_ (.A1(_10948_),
    .A2(_10949_),
    .ZN(_10950_));
 AOI21_X1 _20277_ (.A(_10657_),
    .B1(_10606_),
    .B2(_10564_),
    .ZN(_10951_));
 NAND2_X2 _20278_ (.A1(_10588_),
    .A2(_10660_),
    .ZN(_10952_));
 XNOR2_X1 _20279_ (.A(_10596_),
    .B(_10654_),
    .ZN(_10953_));
 OAI221_X1 _20280_ (.A(_10738_),
    .B1(_10952_),
    .B2(_10564_),
    .C1(_10953_),
    .C2(_10603_),
    .ZN(_10954_));
 AOI221_X1 _20281_ (.A(_10646_),
    .B1(_10950_),
    .B2(_10951_),
    .C1(_10954_),
    .C2(_10695_),
    .ZN(_10955_));
 NOR3_X1 _20282_ (.A1(_10627_),
    .A2(_10947_),
    .A3(_10955_),
    .ZN(_10956_));
 OAI221_X1 _20283_ (.A(_10892_),
    .B1(_10697_),
    .B2(_10632_),
    .C1(_14859_),
    .C2(_10876_),
    .ZN(_10957_));
 AOI21_X1 _20284_ (.A(_10957_),
    .B1(_10635_),
    .B2(_10813_),
    .ZN(_10958_));
 AOI21_X1 _20285_ (.A(_10578_),
    .B1(_10660_),
    .B2(_10452_),
    .ZN(_10959_));
 AOI221_X2 _20286_ (.A(_10596_),
    .B1(_10821_),
    .B2(_10959_),
    .C1(_10622_),
    .C2(_14867_),
    .ZN(_10960_));
 OAI21_X2 _20287_ (.A(_10564_),
    .B1(_10618_),
    .B2(_10619_),
    .ZN(_10961_));
 AOI21_X1 _20288_ (.A(_10570_),
    .B1(_10961_),
    .B2(_10499_),
    .ZN(_10962_));
 OAI21_X1 _20289_ (.A(_10595_),
    .B1(_10629_),
    .B2(_10962_),
    .ZN(_10963_));
 OAI221_X1 _20290_ (.A(_10894_),
    .B1(_10695_),
    .B2(_14864_),
    .C1(_10651_),
    .C2(_10851_),
    .ZN(_10964_));
 OAI221_X1 _20291_ (.A(_10627_),
    .B1(_10960_),
    .B2(_10963_),
    .C1(_10964_),
    .C2(_10728_),
    .ZN(_10965_));
 OAI21_X1 _20292_ (.A(_10511_),
    .B1(_10958_),
    .B2(_10965_),
    .ZN(_10966_));
 NAND2_X1 _20293_ (.A1(_10689_),
    .A2(_10701_),
    .ZN(_10967_));
 AND2_X1 _20294_ (.A1(_10620_),
    .A2(_10821_),
    .ZN(_10968_));
 OAI221_X1 _20295_ (.A(_10948_),
    .B1(_10875_),
    .B2(_10582_),
    .C1(_10968_),
    .C2(_14876_),
    .ZN(_10969_));
 MUX2_X1 _20296_ (.A(_14872_),
    .B(_10747_),
    .S(_10764_),
    .Z(_10970_));
 MUX2_X1 _20297_ (.A(_10969_),
    .B(_10970_),
    .S(_10534_),
    .Z(_10971_));
 OAI221_X1 _20298_ (.A(_10942_),
    .B1(_10956_),
    .B2(_10966_),
    .C1(_10967_),
    .C2(_10971_),
    .ZN(_00052_));
 NOR2_X1 _20299_ (.A1(_10735_),
    .A2(_10585_),
    .ZN(_10972_));
 AOI21_X1 _20300_ (.A(_10972_),
    .B1(_10875_),
    .B2(_14867_),
    .ZN(_10973_));
 NAND2_X1 _20301_ (.A1(_10595_),
    .A2(_10629_),
    .ZN(_10974_));
 OAI21_X1 _20302_ (.A(_10666_),
    .B1(_10973_),
    .B2(_10974_),
    .ZN(_10975_));
 NAND2_X1 _20303_ (.A1(_10532_),
    .A2(_10596_),
    .ZN(_10976_));
 NAND2_X1 _20304_ (.A1(_10564_),
    .A2(_10497_),
    .ZN(_10977_));
 OAI21_X1 _20305_ (.A(_10815_),
    .B1(_10498_),
    .B2(_10602_),
    .ZN(_10978_));
 AOI221_X2 _20306_ (.A(_10976_),
    .B1(_10661_),
    .B2(_10977_),
    .C1(_10978_),
    .C2(_10680_),
    .ZN(_10979_));
 NOR2_X1 _20307_ (.A1(_10609_),
    .A2(_10578_),
    .ZN(_10980_));
 OAI21_X1 _20308_ (.A(_10581_),
    .B1(_10635_),
    .B2(_10980_),
    .ZN(_10981_));
 AOI21_X1 _20309_ (.A(_10797_),
    .B1(_10599_),
    .B2(_10591_),
    .ZN(_10982_));
 NAND2_X1 _20310_ (.A1(_10498_),
    .A2(_10982_),
    .ZN(_10983_));
 AOI21_X1 _20311_ (.A(_10588_),
    .B1(_10691_),
    .B2(_10500_),
    .ZN(_10984_));
 AOI221_X2 _20312_ (.A(_10533_),
    .B1(_10639_),
    .B2(_10981_),
    .C1(_10983_),
    .C2(_10984_),
    .ZN(_10985_));
 NOR3_X1 _20313_ (.A1(_10975_),
    .A2(_10979_),
    .A3(_10985_),
    .ZN(_10986_));
 INV_X1 _20314_ (.A(_10720_),
    .ZN(_10987_));
 AOI21_X1 _20315_ (.A(_10673_),
    .B1(net986),
    .B2(_10599_),
    .ZN(_10988_));
 AOI221_X2 _20316_ (.A(_10729_),
    .B1(_10590_),
    .B2(_10564_),
    .C1(net165),
    .C2(_10660_),
    .ZN(_10989_));
 AOI221_X2 _20317_ (.A(_10645_),
    .B1(_10988_),
    .B2(_10987_),
    .C1(_10989_),
    .C2(_10587_),
    .ZN(_10990_));
 AOI21_X1 _20318_ (.A(_10452_),
    .B1(_10875_),
    .B2(_10952_),
    .ZN(_10991_));
 OAI22_X2 _20319_ (.A1(_10592_),
    .A2(_10851_),
    .B1(_10875_),
    .B2(_14867_),
    .ZN(_10992_));
 NAND3_X1 _20320_ (.A1(net987),
    .A2(_10596_),
    .A3(_10581_),
    .ZN(_10993_));
 MUX2_X1 _20321_ (.A(_10576_),
    .B(_10613_),
    .S(_10546_),
    .Z(_10994_));
 OAI21_X1 _20322_ (.A(_10993_),
    .B1(_10994_),
    .B2(net987),
    .ZN(_10995_));
 AOI221_X2 _20323_ (.A(_10991_),
    .B1(_10992_),
    .B2(_10606_),
    .C1(_14867_),
    .C2(_10995_),
    .ZN(_10996_));
 OAI21_X1 _20324_ (.A(_10990_),
    .B1(_10996_),
    .B2(_10627_),
    .ZN(_10997_));
 MUX2_X1 _20325_ (.A(_10601_),
    .B(_14862_),
    .S(_10580_),
    .Z(_10998_));
 AOI221_X2 _20326_ (.A(_10626_),
    .B1(_10711_),
    .B2(_10450_),
    .C1(_10998_),
    .C2(_10496_),
    .ZN(_10999_));
 OAI21_X1 _20327_ (.A(_10948_),
    .B1(_10724_),
    .B2(_10497_),
    .ZN(_11000_));
 AOI21_X1 _20328_ (.A(_10999_),
    .B1(_11000_),
    .B2(_10626_),
    .ZN(_11001_));
 AOI22_X1 _20329_ (.A1(_10473_),
    .A2(_10563_),
    .B1(_10870_),
    .B2(_10578_),
    .ZN(_11002_));
 MUX2_X1 _20330_ (.A(_10730_),
    .B(_10615_),
    .S(_10576_),
    .Z(_11003_));
 OAI22_X1 _20331_ (.A1(_10602_),
    .A2(_10613_),
    .B1(_11003_),
    .B2(_10578_),
    .ZN(_11004_));
 MUX2_X1 _20332_ (.A(_11002_),
    .B(_11004_),
    .S(_10521_),
    .Z(_11005_));
 AOI221_X2 _20333_ (.A(_10716_),
    .B1(_10894_),
    .B2(_11001_),
    .C1(_11005_),
    .C2(_10892_),
    .ZN(_11006_));
 OAI221_X1 _20334_ (.A(_10595_),
    .B1(_10678_),
    .B2(_10772_),
    .C1(_10880_),
    .C2(_10499_),
    .ZN(_11007_));
 OAI221_X1 _20335_ (.A(_10646_),
    .B1(_10656_),
    .B2(_10678_),
    .C1(_10632_),
    .C2(_10592_),
    .ZN(_11008_));
 AOI21_X1 _20336_ (.A(_10598_),
    .B1(_11007_),
    .B2(_11008_),
    .ZN(_11009_));
 OAI22_X1 _20337_ (.A1(net166),
    .A2(_10851_),
    .B1(_10980_),
    .B2(_10764_),
    .ZN(_11010_));
 AOI21_X1 _20338_ (.A(_10689_),
    .B1(_11010_),
    .B2(_10534_),
    .ZN(_11011_));
 NAND3_X1 _20339_ (.A1(_10623_),
    .A2(_10693_),
    .A3(_10756_),
    .ZN(_11012_));
 NAND3_X1 _20340_ (.A1(_10686_),
    .A2(_10983_),
    .A3(_11012_),
    .ZN(_11013_));
 AOI21_X2 _20341_ (.A(_11009_),
    .B1(_11011_),
    .B2(_11013_),
    .ZN(_11014_));
 AOI221_X2 _20342_ (.A(_10986_),
    .B1(_10997_),
    .B2(_11006_),
    .C1(_11014_),
    .C2(_10701_),
    .ZN(_00053_));
 NOR3_X1 _20343_ (.A1(_14877_),
    .A2(_14886_),
    .A3(_10600_),
    .ZN(_11015_));
 NAND2_X1 _20344_ (.A1(_10586_),
    .A2(_10500_),
    .ZN(_11016_));
 AOI21_X1 _20345_ (.A(_11015_),
    .B1(_11016_),
    .B2(_10721_),
    .ZN(_11017_));
 AND3_X1 _20346_ (.A1(_10631_),
    .A2(_10585_),
    .A3(_10961_),
    .ZN(_11018_));
 MUX2_X1 _20347_ (.A(_10603_),
    .B(_10847_),
    .S(_10680_),
    .Z(_11019_));
 AOI21_X1 _20348_ (.A(_11018_),
    .B1(_11019_),
    .B2(_14883_),
    .ZN(_11020_));
 OAI22_X1 _20349_ (.A1(_10974_),
    .A2(_11017_),
    .B1(_11020_),
    .B2(_10936_),
    .ZN(_11021_));
 OAI21_X1 _20350_ (.A(_10961_),
    .B1(_10660_),
    .B2(_10615_),
    .ZN(_11022_));
 AOI221_X1 _20351_ (.A(_10976_),
    .B1(_11022_),
    .B2(_10500_),
    .C1(_10563_),
    .C2(_10582_),
    .ZN(_11023_));
 OR2_X1 _20352_ (.A1(_10578_),
    .A2(_10690_),
    .ZN(_11024_));
 NOR2_X1 _20353_ (.A1(_10581_),
    .A2(_10671_),
    .ZN(_11025_));
 MUX2_X1 _20354_ (.A(_14874_),
    .B(_10564_),
    .S(_10496_),
    .Z(_11026_));
 AOI221_X1 _20355_ (.A(_10934_),
    .B1(_11024_),
    .B2(_11025_),
    .C1(_11026_),
    .C2(_10607_),
    .ZN(_11027_));
 OR3_X1 _20356_ (.A1(_10628_),
    .A2(_11023_),
    .A3(_11027_),
    .ZN(_11028_));
 OR2_X1 _20357_ (.A1(_11021_),
    .A2(_11028_),
    .ZN(_11029_));
 NOR2_X1 _20358_ (.A1(_10716_),
    .A2(_10627_),
    .ZN(_11030_));
 NOR2_X1 _20359_ (.A1(_10622_),
    .A2(_10570_),
    .ZN(_11031_));
 AOI221_X2 _20360_ (.A(_10597_),
    .B1(_10948_),
    .B2(_11031_),
    .C1(_10896_),
    .C2(_10631_),
    .ZN(_11032_));
 OAI21_X1 _20361_ (.A(_10597_),
    .B1(_10813_),
    .B2(_14879_),
    .ZN(_11033_));
 NOR2_X1 _20362_ (.A1(_10764_),
    .A2(_10917_),
    .ZN(_11034_));
 AOI21_X1 _20363_ (.A(_11033_),
    .B1(_11034_),
    .B2(_10815_),
    .ZN(_11035_));
 NOR3_X1 _20364_ (.A1(_10719_),
    .A2(_11032_),
    .A3(_11035_),
    .ZN(_11036_));
 AOI21_X1 _20365_ (.A(_10498_),
    .B1(_10654_),
    .B2(_10847_),
    .ZN(_11037_));
 AOI22_X2 _20366_ (.A1(_10499_),
    .A2(_10835_),
    .B1(_11037_),
    .B2(_10948_),
    .ZN(_11038_));
 OAI21_X1 _20367_ (.A(_10600_),
    .B1(_10635_),
    .B2(_14859_),
    .ZN(_11039_));
 AOI221_X2 _20368_ (.A(_10595_),
    .B1(_10714_),
    .B2(_11038_),
    .C1(_11039_),
    .C2(_10593_),
    .ZN(_11040_));
 OAI21_X1 _20369_ (.A(_11030_),
    .B1(_11036_),
    .B2(_11040_),
    .ZN(_11041_));
 AOI21_X1 _20370_ (.A(_10623_),
    .B1(_10845_),
    .B2(_10830_),
    .ZN(_11042_));
 OAI21_X1 _20371_ (.A(_10597_),
    .B1(_10614_),
    .B2(_14864_),
    .ZN(_11043_));
 OR2_X1 _20372_ (.A1(_11042_),
    .A2(_11043_),
    .ZN(_11044_));
 NAND3_X1 _20373_ (.A1(_10719_),
    .A2(_10795_),
    .A3(_11044_),
    .ZN(_11045_));
 OAI21_X1 _20374_ (.A(_10879_),
    .B1(_10614_),
    .B2(_10603_),
    .ZN(_11046_));
 AOI22_X1 _20375_ (.A1(_14878_),
    .A2(_10764_),
    .B1(_10661_),
    .B2(_10977_),
    .ZN(_11047_));
 MUX2_X1 _20376_ (.A(_11046_),
    .B(_11047_),
    .S(_10689_),
    .Z(_11048_));
 OAI211_X2 _20377_ (.A(_10701_),
    .B(_11045_),
    .C1(_11048_),
    .C2(_10719_),
    .ZN(_11049_));
 NOR2_X1 _20378_ (.A1(_10521_),
    .A2(_10534_),
    .ZN(_11050_));
 NAND2_X1 _20379_ (.A1(_14859_),
    .A2(_10597_),
    .ZN(_11051_));
 AND3_X1 _20380_ (.A1(_14883_),
    .A2(_10630_),
    .A3(_11051_),
    .ZN(_11052_));
 NAND2_X1 _20381_ (.A1(_10640_),
    .A2(_10588_),
    .ZN(_11053_));
 NOR2_X1 _20382_ (.A1(_10606_),
    .A2(_10788_),
    .ZN(_11054_));
 AOI221_X2 _20383_ (.A(_10657_),
    .B1(_10788_),
    .B2(_11053_),
    .C1(_11054_),
    .C2(_10603_),
    .ZN(_11055_));
 OAI221_X2 _20384_ (.A(_11050_),
    .B1(_11052_),
    .B2(_11055_),
    .C1(_10689_),
    .C2(_10727_),
    .ZN(_11056_));
 NAND3_X1 _20385_ (.A1(_14864_),
    .A2(_14858_),
    .A3(_10629_),
    .ZN(_11057_));
 OAI21_X1 _20386_ (.A(_10623_),
    .B1(_10629_),
    .B2(_10797_),
    .ZN(_11058_));
 OAI221_X2 _20387_ (.A(_11057_),
    .B1(_10952_),
    .B2(_10656_),
    .C1(_14859_),
    .C2(_11058_),
    .ZN(_11059_));
 AOI21_X1 _20388_ (.A(_10683_),
    .B1(_10610_),
    .B2(_14859_),
    .ZN(_11060_));
 OAI221_X1 _20389_ (.A(_10743_),
    .B1(_11060_),
    .B2(net166),
    .C1(_10813_),
    .C2(_10697_),
    .ZN(_11061_));
 AOI22_X1 _20390_ (.A1(_10534_),
    .A2(_11059_),
    .B1(_11061_),
    .B2(_10647_),
    .ZN(_11062_));
 NAND3_X1 _20391_ (.A1(_10666_),
    .A2(_11056_),
    .A3(_11062_),
    .ZN(_11063_));
 NAND4_X1 _20392_ (.A1(_11029_),
    .A2(_11041_),
    .A3(_11049_),
    .A4(_11063_),
    .ZN(_00054_));
 AOI221_X1 _20393_ (.A(_10588_),
    .B1(_10642_),
    .B2(_10615_),
    .C1(_10590_),
    .C2(_14858_),
    .ZN(_11064_));
 OAI21_X1 _20394_ (.A(_10585_),
    .B1(_10851_),
    .B2(_14858_),
    .ZN(_11065_));
 NAND2_X1 _20395_ (.A1(_10668_),
    .A2(_11065_),
    .ZN(_11066_));
 OAI21_X1 _20396_ (.A(_10631_),
    .B1(_10669_),
    .B2(_10797_),
    .ZN(_11067_));
 AOI21_X1 _20397_ (.A(_10606_),
    .B1(_10563_),
    .B2(_10640_),
    .ZN(_11068_));
 AOI221_X1 _20398_ (.A(_10686_),
    .B1(_11064_),
    .B2(_11066_),
    .C1(_11067_),
    .C2(_11068_),
    .ZN(_11069_));
 NAND2_X1 _20399_ (.A1(_10813_),
    .A2(_11026_),
    .ZN(_11070_));
 OAI21_X1 _20400_ (.A(_10764_),
    .B1(_10635_),
    .B2(_10672_),
    .ZN(_11071_));
 NAND3_X1 _20401_ (.A1(_10892_),
    .A2(_11070_),
    .A3(_11071_),
    .ZN(_11072_));
 AOI222_X2 _20402_ (.A1(_10730_),
    .A2(_10642_),
    .B1(_10590_),
    .B2(_14858_),
    .C1(_10876_),
    .C2(_10707_),
    .ZN(_11073_));
 OAI21_X1 _20403_ (.A(_11072_),
    .B1(_11073_),
    .B2(_10936_),
    .ZN(_11074_));
 OAI21_X1 _20404_ (.A(_10666_),
    .B1(_11069_),
    .B2(_11074_),
    .ZN(_11075_));
 INV_X1 _20405_ (.A(_10701_),
    .ZN(_11076_));
 AOI21_X1 _20406_ (.A(_10668_),
    .B1(_10620_),
    .B2(_10650_),
    .ZN(_11077_));
 OAI21_X1 _20407_ (.A(_10629_),
    .B1(_10972_),
    .B2(_11077_),
    .ZN(_11078_));
 OAI21_X1 _20408_ (.A(_10851_),
    .B1(_10656_),
    .B2(_10788_),
    .ZN(_11079_));
 OAI21_X1 _20409_ (.A(_10727_),
    .B1(_10613_),
    .B2(_14867_),
    .ZN(_11080_));
 AOI22_X1 _20410_ (.A1(_14864_),
    .A2(_11079_),
    .B1(_11080_),
    .B2(_10606_),
    .ZN(_11081_));
 AOI21_X1 _20411_ (.A(_10686_),
    .B1(_11078_),
    .B2(_11081_),
    .ZN(_11082_));
 AND4_X1 _20412_ (.A1(_10501_),
    .A2(_10693_),
    .A3(_10844_),
    .A4(_10892_),
    .ZN(_11083_));
 MUX2_X1 _20413_ (.A(_10642_),
    .B(_10590_),
    .S(_10473_),
    .Z(_11084_));
 AOI221_X1 _20414_ (.A(_10936_),
    .B1(_11084_),
    .B2(_10452_),
    .C1(_10711_),
    .C2(_10602_),
    .ZN(_11085_));
 OR4_X2 _20415_ (.A1(_11076_),
    .A2(_11082_),
    .A3(_11083_),
    .A4(_11085_),
    .ZN(_11086_));
 NAND4_X1 _20416_ (.A1(_10582_),
    .A2(_10657_),
    .A3(_10583_),
    .A4(_10584_),
    .ZN(_11087_));
 OAI21_X1 _20417_ (.A(_11087_),
    .B1(_10632_),
    .B2(_14872_),
    .ZN(_11088_));
 AOI21_X1 _20418_ (.A(_10522_),
    .B1(_10653_),
    .B2(_11088_),
    .ZN(_11089_));
 MUX2_X1 _20419_ (.A(net165),
    .B(_10668_),
    .S(_10657_),
    .Z(_11090_));
 OAI221_X1 _20420_ (.A(_10647_),
    .B1(_10678_),
    .B2(_10635_),
    .C1(_11090_),
    .C2(_10813_),
    .ZN(_11091_));
 AND2_X1 _20421_ (.A1(_11089_),
    .A2(_11091_),
    .ZN(_11092_));
 NOR2_X1 _20422_ (.A1(_14886_),
    .A2(_10655_),
    .ZN(_11093_));
 NOR3_X1 _20423_ (.A1(_10600_),
    .A2(_10641_),
    .A3(_10704_),
    .ZN(_11094_));
 NOR3_X1 _20424_ (.A1(_10934_),
    .A2(_11093_),
    .A3(_11094_),
    .ZN(_11095_));
 AOI21_X1 _20425_ (.A(_10723_),
    .B1(_10632_),
    .B2(_14864_),
    .ZN(_11096_));
 OAI21_X1 _20426_ (.A(_10784_),
    .B1(_11096_),
    .B2(_14883_),
    .ZN(_11097_));
 AOI21_X1 _20427_ (.A(_11095_),
    .B1(_11097_),
    .B2(_10894_),
    .ZN(_11098_));
 NOR3_X1 _20428_ (.A1(_14876_),
    .A2(_10570_),
    .A3(_10781_),
    .ZN(_11099_));
 OAI21_X1 _20429_ (.A(_10689_),
    .B1(_10945_),
    .B2(_11099_),
    .ZN(_11100_));
 AOI221_X1 _20430_ (.A(_10589_),
    .B1(_10721_),
    .B2(_11016_),
    .C1(_10607_),
    .C2(_10609_),
    .ZN(_11101_));
 NOR3_X1 _20431_ (.A1(_10534_),
    .A2(_10628_),
    .A3(_11101_),
    .ZN(_11102_));
 AOI22_X2 _20432_ (.A1(_11092_),
    .A2(_11098_),
    .B1(_11100_),
    .B2(_11102_),
    .ZN(_11103_));
 AOI21_X1 _20433_ (.A(_14876_),
    .B1(_10585_),
    .B2(_10961_),
    .ZN(_11104_));
 OAI21_X1 _20434_ (.A(_10705_),
    .B1(_10847_),
    .B2(_10614_),
    .ZN(_11105_));
 OAI21_X1 _20435_ (.A(_10598_),
    .B1(_11104_),
    .B2(_11105_),
    .ZN(_11106_));
 OAI21_X1 _20436_ (.A(_10695_),
    .B1(_10813_),
    .B2(_10591_),
    .ZN(_11107_));
 OAI221_X1 _20437_ (.A(_10689_),
    .B1(_10691_),
    .B2(_11107_),
    .C1(_10757_),
    .C2(_14883_),
    .ZN(_11108_));
 NOR2_X1 _20438_ (.A1(_10719_),
    .A2(_10628_),
    .ZN(_11109_));
 NAND3_X1 _20439_ (.A1(_11106_),
    .A2(_11108_),
    .A3(_11109_),
    .ZN(_11110_));
 AND4_X4 _20440_ (.A1(_11075_),
    .A2(_11086_),
    .A3(_11103_),
    .A4(_11110_),
    .ZN(_00055_));
 INV_X1 _20441_ (.A(_06619_),
    .ZN(_11111_));
 NOR2_X1 _20442_ (.A1(_11111_),
    .A2(_08994_),
    .ZN(_11112_));
 NOR2_X1 _20443_ (.A1(_06619_),
    .A2(_08994_),
    .ZN(_11113_));
 BUF_X4 _20444_ (.A(\sa10_sub[1] ),
    .Z(_11114_));
 BUF_X2 clone102 (.A(_15293_),
    .Z(net102));
 INV_X1 clone65 (.A(net1193),
    .ZN(net65));
 XNOR2_X2 _20447_ (.A(\sa03_sr[0] ),
    .B(\sa10_sub[0] ),
    .ZN(_11117_));
 XNOR2_X2 _20448_ (.A(_11114_),
    .B(_11117_),
    .ZN(_11118_));
 BUF_X8 _20449_ (.A(\sa03_sr[7] ),
    .Z(_11119_));
 BUF_X8 _20450_ (.A(\sa10_sub[7] ),
    .Z(_11120_));
 XNOR2_X2 _20451_ (.A(_11119_),
    .B(_11120_),
    .ZN(_11121_));
 BUF_X4 _20452_ (.A(\sa21_sub[1] ),
    .Z(_11122_));
 XNOR2_X2 _20453_ (.A(_11122_),
    .B(\sa32_sub[1] ),
    .ZN(_11123_));
 XNOR2_X2 _20454_ (.A(_11123_),
    .B(_11121_),
    .ZN(_11124_));
 XNOR2_X2 _20455_ (.A(_11124_),
    .B(_11118_),
    .ZN(_11125_));
 MUX2_X2 _20456_ (.A(_11112_),
    .B(_11113_),
    .S(_11125_),
    .Z(_11126_));
 NAND3_X2 _20457_ (.A1(_06619_),
    .A2(_09728_),
    .A3(_00449_),
    .ZN(_11127_));
 NAND2_X2 _20458_ (.A1(_11111_),
    .A2(_09730_),
    .ZN(_11128_));
 OAI21_X4 _20459_ (.A(_11127_),
    .B1(_11128_),
    .B2(_00449_),
    .ZN(_11129_));
 NOR2_X4 _20460_ (.A1(_11126_),
    .A2(_11129_),
    .ZN(_11130_));
 INV_X8 _20461_ (.A(net883),
    .ZN(_11131_));
 BUF_X2 rebuffer107 (.A(net1211),
    .Z(net590));
 BUF_X16 _20463_ (.A(_11131_),
    .Z(_11133_));
 BUF_X32 _20464_ (.A(_11133_),
    .Z(_11134_));
 BUF_X32 _20465_ (.A(_11134_),
    .Z(_14896_));
 BUF_X4 _20466_ (.A(\sa32_sub[0] ),
    .Z(_11135_));
 BUF_X4 _20467_ (.A(\sa21_sub[0] ),
    .Z(_11136_));
 XNOR2_X2 _20468_ (.A(_11136_),
    .B(\sa10_sub[0] ),
    .ZN(_11137_));
 XNOR2_X1 _20469_ (.A(_11135_),
    .B(net966),
    .ZN(_11138_));
 XOR2_X2 _20470_ (.A(_11119_),
    .B(_11120_),
    .Z(_11139_));
 NAND3_X1 _20471_ (.A1(net786),
    .A2(_09023_),
    .A3(_11139_),
    .ZN(_11140_));
 NOR2_X1 _20472_ (.A1(net787),
    .A2(_09027_),
    .ZN(_11141_));
 NAND2_X1 _20473_ (.A1(net577),
    .A2(_11141_),
    .ZN(_11142_));
 AOI21_X1 _20474_ (.A(_11138_),
    .B1(_11140_),
    .B2(_11142_),
    .ZN(_11143_));
 XOR2_X2 _20475_ (.A(net579),
    .B(_11136_),
    .Z(_11144_));
 XNOR2_X1 _20476_ (.A(_11135_),
    .B(_11144_),
    .ZN(_11145_));
 NAND2_X1 _20477_ (.A1(_11139_),
    .A2(_11141_),
    .ZN(_11146_));
 NAND3_X1 _20478_ (.A1(net795),
    .A2(_09074_),
    .A3(net576),
    .ZN(_11147_));
 AOI21_X1 _20479_ (.A(_11145_),
    .B1(_11146_),
    .B2(_11147_),
    .ZN(_11148_));
 INV_X1 _20480_ (.A(\u0.tmp_w[24] ),
    .ZN(_11149_));
 NAND3_X1 _20481_ (.A1(_11149_),
    .A2(_08973_),
    .A3(_00450_),
    .ZN(_11150_));
 NAND2_X1 _20482_ (.A1(\u0.tmp_w[24] ),
    .A2(_09727_),
    .ZN(_11151_));
 OAI21_X1 _20483_ (.A(_11150_),
    .B1(_11151_),
    .B2(_00450_),
    .ZN(_11152_));
 OR3_X2 _20484_ (.A1(_11143_),
    .A2(_11148_),
    .A3(_11152_),
    .ZN(_11153_));
 INV_X2 _20485_ (.A(_11153_),
    .ZN(_11154_));
 BUF_X8 _20486_ (.A(_11154_),
    .Z(_11155_));
 BUF_X4 _20487_ (.A(_11155_),
    .Z(_14899_));
 INV_X2 _20488_ (.A(_06635_),
    .ZN(_11156_));
 NOR3_X1 _20489_ (.A1(_11156_),
    .A2(_09099_),
    .A3(_00451_),
    .ZN(_11157_));
 BUF_X4 _20490_ (.A(\sa10_sub[2] ),
    .Z(_11158_));
 BUF_X4 _20491_ (.A(\sa21_sub[2] ),
    .Z(_11159_));
 XNOR2_X2 _20492_ (.A(_11158_),
    .B(_11159_),
    .ZN(_11160_));
 NOR3_X1 _20493_ (.A1(_11156_),
    .A2(_08992_),
    .A3(_11160_),
    .ZN(_11161_));
 XOR2_X2 _20494_ (.A(_11158_),
    .B(_11159_),
    .Z(_11162_));
 NOR3_X1 _20495_ (.A1(_11156_),
    .A2(_08992_),
    .A3(_11162_),
    .ZN(_11163_));
 CLKBUF_X3 _20496_ (.A(\sa32_sub[2] ),
    .Z(_11164_));
 BUF_X1 rebuffer191 (.A(\sa03_sr[1] ),
    .Z(net657));
 XNOR2_X2 _20498_ (.A(\sa03_sr[1] ),
    .B(_11114_),
    .ZN(_11166_));
 XNOR2_X2 _20499_ (.A(_11164_),
    .B(net660),
    .ZN(_11167_));
 MUX2_X1 _20500_ (.A(_11161_),
    .B(_11163_),
    .S(_11167_),
    .Z(_11168_));
 NAND2_X1 _20501_ (.A1(_09022_),
    .A2(_11162_),
    .ZN(_11169_));
 NAND2_X1 _20502_ (.A1(_09022_),
    .A2(_11160_),
    .ZN(_11170_));
 MUX2_X1 _20503_ (.A(_11169_),
    .B(_11170_),
    .S(_11167_),
    .Z(_11171_));
 NOR2_X1 _20504_ (.A1(_09099_),
    .A2(_00451_),
    .ZN(_11172_));
 NOR2_X1 _20505_ (.A1(_06635_),
    .A2(_11172_),
    .ZN(_11173_));
 AOI211_X2 _20506_ (.A(_11157_),
    .B(_11168_),
    .C1(_11171_),
    .C2(_11173_),
    .ZN(_11174_));
 INV_X2 _20507_ (.A(_11174_),
    .ZN(_11175_));
 BUF_X4 _20508_ (.A(_11175_),
    .Z(_11176_));
 CLKBUF_X3 _20509_ (.A(_11176_),
    .Z(_11177_));
 CLKBUF_X3 _20510_ (.A(_11177_),
    .Z(_11178_));
 BUF_X4 _20511_ (.A(_11178_),
    .Z(_14915_));
 BUF_X8 _20512_ (.A(_11153_),
    .Z(_11179_));
 BUF_X4 _20513_ (.A(_11179_),
    .Z(_14890_));
 BUF_X4 _20514_ (.A(_11174_),
    .Z(_11180_));
 BUF_X4 _20515_ (.A(_11180_),
    .Z(_11181_));
 BUF_X4 _20516_ (.A(_11181_),
    .Z(_11182_));
 BUF_X4 _20517_ (.A(_11182_),
    .Z(_14908_));
 BUF_X8 _20518_ (.A(\sa21_sub[7] ),
    .Z(_11183_));
 BUF_X8 _20519_ (.A(\sa32_sub[7] ),
    .Z(_11184_));
 XNOR2_X2 _20520_ (.A(_11183_),
    .B(_11184_),
    .ZN(_11185_));
 CLKBUF_X3 _20521_ (.A(\sa10_sub[6] ),
    .Z(_11186_));
 BUF_X2 _20522_ (.A(\sa03_sr[6] ),
    .Z(_11187_));
 XNOR2_X1 _20523_ (.A(_11186_),
    .B(_11187_),
    .ZN(_11188_));
 XNOR2_X1 _20524_ (.A(_11185_),
    .B(_11188_),
    .ZN(_11189_));
 XNOR2_X1 _20525_ (.A(_11120_),
    .B(_11189_),
    .ZN(_11190_));
 BUF_X32 _20526_ (.A(_09856_),
    .Z(_11191_));
 BUF_X4 _20527_ (.A(_11191_),
    .Z(_11192_));
 MUX2_X2 _20528_ (.A(\text_in_r[31] ),
    .B(_11190_),
    .S(_11192_),
    .Z(_11193_));
 XOR2_X2 _20529_ (.A(_06708_),
    .B(_11193_),
    .Z(_11194_));
 INV_X1 _20530_ (.A(_06699_),
    .ZN(_11195_));
 NOR2_X1 _20531_ (.A1(_11195_),
    .A2(_09136_),
    .ZN(_11196_));
 NOR2_X1 _20532_ (.A1(_06699_),
    .A2(_09136_),
    .ZN(_11197_));
 BUF_X4 _20533_ (.A(\sa32_sub[6] ),
    .Z(_11198_));
 BUF_X2 _20534_ (.A(\sa21_sub[6] ),
    .Z(_11199_));
 XNOR2_X2 _20535_ (.A(_11186_),
    .B(_11199_),
    .ZN(_11200_));
 CLKBUF_X3 _20536_ (.A(\sa10_sub[5] ),
    .Z(_11201_));
 CLKBUF_X3 _20537_ (.A(\sa03_sr[5] ),
    .Z(_11202_));
 XNOR2_X2 _20538_ (.A(_11201_),
    .B(_11202_),
    .ZN(_11203_));
 XNOR2_X1 _20539_ (.A(_11200_),
    .B(_11203_),
    .ZN(_11204_));
 XNOR2_X1 _20540_ (.A(_11198_),
    .B(_11204_),
    .ZN(_11205_));
 MUX2_X2 _20541_ (.A(_11196_),
    .B(_11197_),
    .S(_11205_),
    .Z(_11206_));
 BUF_X4 _20542_ (.A(_11192_),
    .Z(_11207_));
 NOR3_X4 _20543_ (.A1(_11195_),
    .A2(_11207_),
    .A3(\text_in_r[30] ),
    .ZN(_11208_));
 AND3_X1 _20544_ (.A1(_11195_),
    .A2(_09136_),
    .A3(\text_in_r[30] ),
    .ZN(_11209_));
 NOR3_X4 _20545_ (.A1(_11206_),
    .A2(_11208_),
    .A3(_11209_),
    .ZN(_11210_));
 NOR2_X2 _20546_ (.A1(_11194_),
    .A2(_11210_),
    .ZN(_11211_));
 INV_X1 _20547_ (.A(_11211_),
    .ZN(_11212_));
 BUF_X8 clone49 (.A(net829),
    .Z(net49));
 BUF_X4 _20549_ (.A(_14897_),
    .Z(_11214_));
 BUF_X4 _20550_ (.A(_11180_),
    .Z(_11215_));
 NOR2_X1 _20551_ (.A1(_06654_),
    .A2(_08993_),
    .ZN(_11216_));
 INV_X1 _20552_ (.A(_06654_),
    .ZN(_11217_));
 NOR2_X1 _20553_ (.A1(_11217_),
    .A2(_08993_),
    .ZN(_11218_));
 BUF_X4 _20554_ (.A(\sa03_sr[2] ),
    .Z(_11219_));
 BUF_X2 _20555_ (.A(\sa21_sub[3] ),
    .Z(_11220_));
 XNOR2_X1 _20556_ (.A(_11219_),
    .B(_11220_),
    .ZN(_11221_));
 XNOR2_X2 _20557_ (.A(_11119_),
    .B(_11221_),
    .ZN(_11222_));
 CLKBUF_X3 _20558_ (.A(\sa10_sub[3] ),
    .Z(_11223_));
 XOR2_X2 _20559_ (.A(_11120_),
    .B(_11223_),
    .Z(_11224_));
 BUF_X2 _20560_ (.A(\sa32_sub[3] ),
    .Z(_11225_));
 XNOR2_X1 _20561_ (.A(_11158_),
    .B(_11225_),
    .ZN(_11226_));
 XNOR2_X1 _20562_ (.A(_11224_),
    .B(_11226_),
    .ZN(_11227_));
 XNOR2_X1 _20563_ (.A(_11222_),
    .B(_11227_),
    .ZN(_11228_));
 MUX2_X1 _20564_ (.A(_11216_),
    .B(_11218_),
    .S(_11228_),
    .Z(_11229_));
 BUF_X8 _20565_ (.A(_11229_),
    .Z(_11230_));
 BUF_X8 _20566_ (.A(_11230_),
    .Z(_11231_));
 OR3_X2 _20567_ (.A1(_11217_),
    .A2(_09099_),
    .A3(\text_in_r[27] ),
    .ZN(_11232_));
 NAND3_X2 _20568_ (.A1(_11217_),
    .A2(_09102_),
    .A3(\text_in_r[27] ),
    .ZN(_11233_));
 NAND2_X4 _20569_ (.A1(_11232_),
    .A2(_11233_),
    .ZN(_11234_));
 BUF_X8 _20570_ (.A(_11234_),
    .Z(_11235_));
 OAI21_X4 _20571_ (.A(_11215_),
    .B1(_11231_),
    .B2(_11235_),
    .ZN(_11236_));
 BUF_X4 _20572_ (.A(_11176_),
    .Z(_11237_));
 NAND2_X1 _20573_ (.A1(_14890_),
    .A2(_11237_),
    .ZN(_11238_));
 NOR2_X4 _20574_ (.A1(_11230_),
    .A2(_11234_),
    .ZN(_11239_));
 NOR2_X2 _20575_ (.A1(net649),
    .A2(_11239_),
    .ZN(_11240_));
 OAI22_X1 _20576_ (.A1(_11214_),
    .A2(_11236_),
    .B1(_11238_),
    .B2(_11240_),
    .ZN(_11241_));
 INV_X1 _20577_ (.A(_06670_),
    .ZN(_11242_));
 NAND2_X1 _20578_ (.A1(_11242_),
    .A2(_11192_),
    .ZN(_11243_));
 NAND2_X1 _20579_ (.A1(_06670_),
    .A2(_11192_),
    .ZN(_11244_));
 BUF_X2 _20580_ (.A(\sa03_sr[3] ),
    .Z(_11245_));
 BUF_X4 _20581_ (.A(\sa21_sub[4] ),
    .Z(_11246_));
 XNOR2_X1 _20582_ (.A(_11245_),
    .B(_11246_),
    .ZN(_11247_));
 XNOR2_X2 _20583_ (.A(_11119_),
    .B(_11247_),
    .ZN(_11248_));
 CLKBUF_X3 _20584_ (.A(\sa10_sub[4] ),
    .Z(_11249_));
 BUF_X4 _20585_ (.A(\sa32_sub[4] ),
    .Z(_11250_));
 XNOR2_X1 _20586_ (.A(_11249_),
    .B(_11250_),
    .ZN(_11251_));
 XNOR2_X2 _20587_ (.A(_11224_),
    .B(_11251_),
    .ZN(_11252_));
 XNOR2_X2 _20588_ (.A(_11248_),
    .B(_11252_),
    .ZN(_11253_));
 MUX2_X2 _20589_ (.A(_11243_),
    .B(_11244_),
    .S(_11253_),
    .Z(_11254_));
 NAND3_X2 _20590_ (.A1(_11242_),
    .A2(_09135_),
    .A3(\text_in_r[28] ),
    .ZN(_11255_));
 NAND2_X1 _20591_ (.A1(_06670_),
    .A2(net582),
    .ZN(_11256_));
 OAI21_X4 _20592_ (.A(_11255_),
    .B1(_11256_),
    .B2(\text_in_r[28] ),
    .ZN(_11257_));
 INV_X2 _20593_ (.A(_11257_),
    .ZN(_11258_));
 NAND2_X4 _20594_ (.A1(_11254_),
    .A2(_11258_),
    .ZN(_11259_));
 AND2_X1 _20595_ (.A1(_08974_),
    .A2(\text_in_r[29] ),
    .ZN(_11260_));
 CLKBUF_X3 _20596_ (.A(\sa21_sub[5] ),
    .Z(_11261_));
 BUF_X4 _20597_ (.A(\sa32_sub[5] ),
    .Z(_11262_));
 XNOR2_X2 _20598_ (.A(_11261_),
    .B(_11262_),
    .ZN(_11263_));
 XNOR2_X2 _20599_ (.A(_11249_),
    .B(_11263_),
    .ZN(_11264_));
 CLKBUF_X3 _20600_ (.A(\sa03_sr[4] ),
    .Z(_11265_));
 XNOR2_X1 _20601_ (.A(_11265_),
    .B(_11201_),
    .ZN(_11266_));
 XNOR2_X2 _20602_ (.A(_11264_),
    .B(_11266_),
    .ZN(_11267_));
 AOI21_X4 _20603_ (.A(_11260_),
    .B1(_11267_),
    .B2(_09076_),
    .ZN(_11268_));
 XOR2_X2 _20604_ (.A(_06685_),
    .B(_11268_),
    .Z(_11269_));
 NOR2_X2 _20605_ (.A1(_11259_),
    .A2(_11269_),
    .ZN(_11270_));
 AOI21_X1 _20606_ (.A(_11212_),
    .B1(_11241_),
    .B2(_11270_),
    .ZN(_11271_));
 NOR2_X1 _20607_ (.A1(_11154_),
    .A2(_11180_),
    .ZN(_11272_));
 AND2_X1 _20608_ (.A1(_11232_),
    .A2(_11233_),
    .ZN(_11273_));
 BUF_X4 _20609_ (.A(_11273_),
    .Z(_11274_));
 NAND2_X1 _20610_ (.A1(_11217_),
    .A2(_09195_),
    .ZN(_11275_));
 NAND2_X1 _20611_ (.A1(_06654_),
    .A2(_09195_),
    .ZN(_11276_));
 MUX2_X1 _20612_ (.A(_11275_),
    .B(_11276_),
    .S(_11228_),
    .Z(_11277_));
 BUF_X4 _20613_ (.A(_11277_),
    .Z(_11278_));
 NOR2_X4 _20614_ (.A1(_11179_),
    .A2(_11175_),
    .ZN(_11279_));
 AOI221_X2 _20615_ (.A(_11272_),
    .B1(_11274_),
    .B2(_11278_),
    .C1(_11131_),
    .C2(_11279_),
    .ZN(_11280_));
 NOR2_X2 _20616_ (.A1(_11259_),
    .A2(_11280_),
    .ZN(_11281_));
 NAND2_X1 _20617_ (.A1(net649),
    .A2(_11176_),
    .ZN(_11282_));
 BUF_X4 _20618_ (.A(_14894_),
    .Z(_11283_));
 OAI21_X1 _20619_ (.A(_11282_),
    .B1(_14915_),
    .B2(_11283_),
    .ZN(_11284_));
 NAND2_X4 _20620_ (.A1(_11278_),
    .A2(_11274_),
    .ZN(_11285_));
 BUF_X4 _20621_ (.A(_11285_),
    .Z(_11286_));
 CLKBUF_X3 _20622_ (.A(_11286_),
    .Z(_11287_));
 OAI21_X1 _20623_ (.A(_11281_),
    .B1(_11284_),
    .B2(_11287_),
    .ZN(_11288_));
 XNOR2_X2 _20624_ (.A(_06685_),
    .B(_11268_),
    .ZN(_11289_));
 BUF_X4 _20625_ (.A(_11289_),
    .Z(_11290_));
 BUF_X4 _20626_ (.A(_11290_),
    .Z(_11291_));
 CLKBUF_X3 _20627_ (.A(_11291_),
    .Z(_11292_));
 NOR2_X1 _20628_ (.A1(_06670_),
    .A2(_08996_),
    .ZN(_11293_));
 NOR2_X1 _20629_ (.A1(_11242_),
    .A2(_08996_),
    .ZN(_11294_));
 MUX2_X2 _20630_ (.A(_11293_),
    .B(_11294_),
    .S(_11253_),
    .Z(_11295_));
 NOR2_X4 _20631_ (.A1(_11295_),
    .A2(_11257_),
    .ZN(_11296_));
 BUF_X4 _20632_ (.A(_11296_),
    .Z(_11297_));
 CLKBUF_X3 _20633_ (.A(_11297_),
    .Z(_11298_));
 BUF_X4 _20634_ (.A(_11269_),
    .Z(_11299_));
 CLKBUF_X3 _20635_ (.A(_11299_),
    .Z(_11300_));
 NOR2_X1 _20636_ (.A1(_14896_),
    .A2(_11287_),
    .ZN(_11301_));
 TAPCELL_X1 PHY_EDGE_ROW_2_Right_2 ();
 BUF_X4 _20638_ (.A(_11239_),
    .Z(_11303_));
 BUF_X4 _20639_ (.A(_11303_),
    .Z(_11304_));
 MUX2_X1 _20640_ (.A(net562),
    .B(_14896_),
    .S(_11304_),
    .Z(_11305_));
 OAI221_X1 _20641_ (.A(_11300_),
    .B1(_11301_),
    .B2(_11238_),
    .C1(_11305_),
    .C2(_14915_),
    .ZN(_11306_));
 NOR3_X4 _20642_ (.A1(_11179_),
    .A2(_11230_),
    .A3(_11234_),
    .ZN(_11307_));
 BUF_X8 _20643_ (.A(_11130_),
    .Z(_11308_));
 MUX2_X1 _20644_ (.A(_14906_),
    .B(net162),
    .S(_11303_),
    .Z(_11309_));
 AOI21_X4 _20645_ (.A(_11176_),
    .B1(_11278_),
    .B2(_11274_),
    .ZN(_11310_));
 INV_X2 clone43 (.A(_14661_),
    .ZN(net43));
 BUF_X8 _20647_ (.A(net10),
    .Z(_11312_));
 AOI221_X2 _20648_ (.A(_11307_),
    .B1(_11309_),
    .B2(_11178_),
    .C1(_11310_),
    .C2(net734),
    .ZN(_11313_));
 OAI21_X2 _20649_ (.A(_11306_),
    .B1(_11300_),
    .B2(_11313_),
    .ZN(_11314_));
 OAI221_X2 _20650_ (.A(_11271_),
    .B1(_11288_),
    .B2(_11292_),
    .C1(_11314_),
    .C2(_11298_),
    .ZN(_11315_));
 CLKBUF_X3 _20651_ (.A(_11210_),
    .Z(_11316_));
 BUF_X4 _20652_ (.A(_11269_),
    .Z(_11317_));
 CLKBUF_X3 _20653_ (.A(_11317_),
    .Z(_11318_));
 BUF_X4 _20654_ (.A(_11259_),
    .Z(_11319_));
 NAND3_X1 _20655_ (.A1(_14913_),
    .A2(_11319_),
    .A3(_11287_),
    .ZN(_11320_));
 NAND3_X1 _20656_ (.A1(_11316_),
    .A2(_11318_),
    .A3(_11320_),
    .ZN(_11321_));
 BUF_X4 _20657_ (.A(_14892_),
    .Z(_11322_));
 OAI21_X4 _20658_ (.A(_11155_),
    .B1(_11231_),
    .B2(_11235_),
    .ZN(_11323_));
 NAND3_X2 _20659_ (.A1(_11283_),
    .A2(_11278_),
    .A3(_11274_),
    .ZN(_11324_));
 AND2_X1 _20660_ (.A1(_11323_),
    .A2(_11324_),
    .ZN(_11325_));
 BUF_X4 _20661_ (.A(_11215_),
    .Z(_11326_));
 BUF_X4 _20662_ (.A(_11326_),
    .Z(_11327_));
 OAI22_X2 _20663_ (.A1(_11322_),
    .A2(_11236_),
    .B1(_11325_),
    .B2(_11327_),
    .ZN(_11328_));
 BUF_X4 _20664_ (.A(_11297_),
    .Z(_11329_));
 BUF_X4 _20665_ (.A(_11304_),
    .Z(_11330_));
 BUF_X4 _20666_ (.A(_11176_),
    .Z(_11331_));
 BUF_X4 _20667_ (.A(_11331_),
    .Z(_11332_));
 BUF_X4 _20668_ (.A(_11332_),
    .Z(_11333_));
 MUX2_X1 _20669_ (.A(net734),
    .B(_11214_),
    .S(_11296_),
    .Z(_11334_));
 NAND2_X1 _20670_ (.A1(net651),
    .A2(_14890_),
    .ZN(_11335_));
 CLKBUF_X3 _20671_ (.A(_11259_),
    .Z(_11336_));
 NOR2_X1 _20672_ (.A1(_11177_),
    .A2(_11336_),
    .ZN(_11337_));
 AOI22_X1 _20673_ (.A1(_11333_),
    .A2(_11334_),
    .B1(_11335_),
    .B2(_11337_),
    .ZN(_11338_));
 INV_X1 _20674_ (.A(_11338_),
    .ZN(_11339_));
 AOI221_X2 _20675_ (.A(_11321_),
    .B1(_11328_),
    .B2(_11329_),
    .C1(_11330_),
    .C2(_11339_),
    .ZN(_11340_));
 CLKBUF_X3 _20676_ (.A(_14900_),
    .Z(_11341_));
 INV_X1 _20677_ (.A(_11341_),
    .ZN(_11342_));
 OAI21_X2 _20678_ (.A(_11342_),
    .B1(_11231_),
    .B2(_11235_),
    .ZN(_11343_));
 NOR3_X4 _20679_ (.A1(net648),
    .A2(_11230_),
    .A3(_11234_),
    .ZN(_11344_));
 NOR2_X2 _20680_ (.A1(_11344_),
    .A2(_11180_),
    .ZN(_11345_));
 BUF_X4 _20681_ (.A(_11278_),
    .Z(_11346_));
 BUF_X4 _20682_ (.A(_11274_),
    .Z(_11347_));
 AOI21_X2 _20683_ (.A(_11179_),
    .B1(_11346_),
    .B2(_11347_),
    .ZN(_11348_));
 AOI21_X1 _20684_ (.A(_11348_),
    .B1(_11303_),
    .B2(net162),
    .ZN(_11349_));
 AOI221_X1 _20685_ (.A(_11259_),
    .B1(_11343_),
    .B2(_11345_),
    .C1(_11349_),
    .C2(_11326_),
    .ZN(_11350_));
 OAI21_X4 _20686_ (.A(net852),
    .B1(_11230_),
    .B2(_11234_),
    .ZN(_11351_));
 AND2_X4 _20687_ (.A1(_11180_),
    .A2(_11351_),
    .ZN(_11352_));
 NOR3_X2 _20688_ (.A1(_11180_),
    .A2(_11230_),
    .A3(_11234_),
    .ZN(_11353_));
 CLKBUF_X3 _20689_ (.A(_11353_),
    .Z(_11354_));
 AOI221_X2 _20690_ (.A(_11296_),
    .B1(_11324_),
    .B2(_11352_),
    .C1(_11354_),
    .C2(_11322_),
    .ZN(_11355_));
 OR4_X2 _20691_ (.A1(_11350_),
    .A2(_11355_),
    .A3(_11316_),
    .A4(_11318_),
    .ZN(_11356_));
 OR3_X4 _20692_ (.A1(_11206_),
    .A2(_11208_),
    .A3(_11209_),
    .ZN(_11357_));
 CLKBUF_X3 _20693_ (.A(_11357_),
    .Z(_11358_));
 NAND2_X1 _20694_ (.A1(_11358_),
    .A2(_11299_),
    .ZN(_11359_));
 AOI21_X2 _20695_ (.A(_11154_),
    .B1(_11278_),
    .B2(_11274_),
    .ZN(_11360_));
 BUF_X4 _20696_ (.A(_11360_),
    .Z(_11361_));
 NAND2_X1 _20697_ (.A1(_11296_),
    .A2(_11361_),
    .ZN(_11362_));
 NOR3_X4 _20698_ (.A1(net851),
    .A2(_11230_),
    .A3(_11234_),
    .ZN(_11363_));
 NOR2_X1 _20699_ (.A1(_14908_),
    .A2(_11363_),
    .ZN(_11364_));
 AOI21_X1 _20700_ (.A(_11359_),
    .B1(_11362_),
    .B2(_11364_),
    .ZN(_11365_));
 OAI21_X4 _20701_ (.A(net10),
    .B1(_11231_),
    .B2(_11235_),
    .ZN(_11366_));
 BUF_X2 _20702_ (.A(_14902_),
    .Z(_11367_));
 BUF_X4 _20703_ (.A(_11367_),
    .Z(_11368_));
 NAND3_X2 _20704_ (.A1(_11368_),
    .A2(_11346_),
    .A3(_11347_),
    .ZN(_11369_));
 AOI21_X1 _20705_ (.A(_11333_),
    .B1(net733),
    .B2(_11369_),
    .ZN(_11370_));
 NOR2_X1 _20706_ (.A1(_11298_),
    .A2(_11370_),
    .ZN(_11371_));
 OAI21_X1 _20707_ (.A(_11365_),
    .B1(_11371_),
    .B2(_11281_),
    .ZN(_11372_));
 BUF_X4 _20708_ (.A(_11285_),
    .Z(_11373_));
 CLKBUF_X3 _20709_ (.A(_11373_),
    .Z(_11374_));
 OAI21_X4 _20710_ (.A(_11179_),
    .B1(_11231_),
    .B2(_11235_),
    .ZN(_11375_));
 BUF_X16 _20711_ (.A(_11308_),
    .Z(_11376_));
 OAI221_X1 _20712_ (.A(_11327_),
    .B1(_11374_),
    .B2(_11283_),
    .C1(_11375_),
    .C2(_11376_),
    .ZN(_11377_));
 AOI21_X4 _20713_ (.A(_11180_),
    .B1(_11278_),
    .B2(_11274_),
    .ZN(_11378_));
 NAND2_X1 _20714_ (.A1(_11368_),
    .A2(_11378_),
    .ZN(_11379_));
 NAND4_X1 _20715_ (.A1(_11316_),
    .A2(_11270_),
    .A3(_11377_),
    .A4(_11379_),
    .ZN(_11380_));
 NAND2_X1 _20716_ (.A1(_11342_),
    .A2(_11354_),
    .ZN(_11381_));
 NAND3_X4 _20717_ (.A1(_11179_),
    .A2(_11346_),
    .A3(_11347_),
    .ZN(_11382_));
 OAI221_X2 _20718_ (.A(_11327_),
    .B1(_11304_),
    .B2(_11283_),
    .C1(_11382_),
    .C2(_11376_),
    .ZN(_11383_));
 NOR2_X1 _20719_ (.A1(_11297_),
    .A2(_11299_),
    .ZN(_11384_));
 NAND4_X1 _20720_ (.A1(_11316_),
    .A2(_11381_),
    .A3(_11383_),
    .A4(_11384_),
    .ZN(_11385_));
 AND3_X1 _20721_ (.A1(_11194_),
    .A2(_11380_),
    .A3(_11385_),
    .ZN(_11386_));
 NAND3_X2 _20722_ (.A1(_11356_),
    .A2(_11372_),
    .A3(_11386_),
    .ZN(_11387_));
 XNOR2_X2 _20723_ (.A(_06708_),
    .B(_11193_),
    .ZN(_11388_));
 NAND2_X1 _20724_ (.A1(_11388_),
    .A2(_11316_),
    .ZN(_11389_));
 BUF_X4 _20725_ (.A(_11296_),
    .Z(_11390_));
 CLKBUF_X3 _20726_ (.A(_11289_),
    .Z(_11391_));
 NAND2_X1 _20727_ (.A1(_11390_),
    .A2(_11391_),
    .ZN(_11392_));
 NOR2_X1 _20728_ (.A1(_11332_),
    .A2(_11344_),
    .ZN(_11393_));
 OAI21_X1 _20729_ (.A(_11341_),
    .B1(_11231_),
    .B2(_11235_),
    .ZN(_11394_));
 NAND2_X1 _20730_ (.A1(_11393_),
    .A2(_11394_),
    .ZN(_11395_));
 NAND2_X2 _20731_ (.A1(_11131_),
    .A2(_11307_),
    .ZN(_11396_));
 NAND2_X2 _20732_ (.A1(_11322_),
    .A2(_11373_),
    .ZN(_11397_));
 NAND3_X1 _20733_ (.A1(_11333_),
    .A2(_11396_),
    .A3(_11397_),
    .ZN(_11398_));
 AOI21_X1 _20734_ (.A(_11392_),
    .B1(_11395_),
    .B2(_11398_),
    .ZN(_11399_));
 NOR3_X4 _20735_ (.A1(_11175_),
    .A2(_11230_),
    .A3(_11234_),
    .ZN(_11400_));
 NOR2_X4 _20736_ (.A1(_11378_),
    .A2(_11400_),
    .ZN(_11401_));
 INV_X8 _20737_ (.A(net10),
    .ZN(_11402_));
 OAI221_X2 _20738_ (.A(_11381_),
    .B1(_11401_),
    .B2(_11322_),
    .C1(_11236_),
    .C2(net161),
    .ZN(_11403_));
 NOR2_X2 _20739_ (.A1(_11319_),
    .A2(_11290_),
    .ZN(_11404_));
 CLKBUF_X3 _20740_ (.A(_11319_),
    .Z(_11405_));
 BUF_X4 _20741_ (.A(_11181_),
    .Z(_11406_));
 OAI21_X1 _20742_ (.A(_11406_),
    .B1(_11317_),
    .B2(_14899_),
    .ZN(_11407_));
 NOR2_X2 _20743_ (.A1(_11179_),
    .A2(_11215_),
    .ZN(_11408_));
 NOR2_X2 _20744_ (.A1(_11331_),
    .A2(_11289_),
    .ZN(_11409_));
 AOI222_X2 _20745_ (.A1(_11134_),
    .A2(_11407_),
    .B1(_11408_),
    .B2(_11391_),
    .C1(_11409_),
    .C2(net734),
    .ZN(_11410_));
 NOR2_X1 _20746_ (.A1(net649),
    .A2(_11155_),
    .ZN(_11411_));
 OAI21_X1 _20747_ (.A(_11290_),
    .B1(_11279_),
    .B2(_11411_),
    .ZN(_11412_));
 CLKBUF_X3 _20748_ (.A(_11239_),
    .Z(_11413_));
 CLKBUF_X3 _20749_ (.A(_11413_),
    .Z(_11414_));
 NOR3_X1 _20750_ (.A1(_11312_),
    .A2(_11406_),
    .A3(_11391_),
    .ZN(_11415_));
 NOR2_X1 _20751_ (.A1(_11414_),
    .A2(_11415_),
    .ZN(_11416_));
 AOI22_X2 _20752_ (.A1(_11330_),
    .A2(_11410_),
    .B1(_11412_),
    .B2(_11416_),
    .ZN(_11417_));
 AOI221_X2 _20753_ (.A(_11399_),
    .B1(_11403_),
    .B2(_11404_),
    .C1(_11405_),
    .C2(_11417_),
    .ZN(_11418_));
 OAI221_X2 _20754_ (.A(_11315_),
    .B1(_11340_),
    .B2(_11387_),
    .C1(_11389_),
    .C2(_11418_),
    .ZN(_00056_));
 NOR2_X2 _20755_ (.A1(_11388_),
    .A2(_11357_),
    .ZN(_11419_));
 BUF_X4 _20756_ (.A(_11130_),
    .Z(_11420_));
 AOI21_X1 _20757_ (.A(_11420_),
    .B1(_11177_),
    .B2(_11375_),
    .ZN(_11421_));
 OAI221_X1 _20758_ (.A(_11270_),
    .B1(_11382_),
    .B2(net651),
    .C1(_11237_),
    .C2(_11413_),
    .ZN(_11422_));
 OAI21_X1 _20759_ (.A(_11419_),
    .B1(_11421_),
    .B2(_11422_),
    .ZN(_11423_));
 NAND3_X2 _20760_ (.A1(_14897_),
    .A2(_11346_),
    .A3(_11347_),
    .ZN(_11424_));
 AOI21_X1 _20761_ (.A(_11331_),
    .B1(_11366_),
    .B2(_11424_),
    .ZN(_11425_));
 NOR3_X1 _20762_ (.A1(_11181_),
    .A2(_11307_),
    .A3(_11361_),
    .ZN(_11426_));
 OAI21_X1 _20763_ (.A(_11391_),
    .B1(_11425_),
    .B2(_11426_),
    .ZN(_11427_));
 NAND2_X1 _20764_ (.A1(_11331_),
    .A2(_11303_),
    .ZN(_11428_));
 OAI22_X1 _20765_ (.A1(_11214_),
    .A2(_11428_),
    .B1(_11401_),
    .B2(_11420_),
    .ZN(_11429_));
 OAI21_X1 _20766_ (.A(_11427_),
    .B1(_11429_),
    .B2(_11290_),
    .ZN(_11430_));
 AOI21_X2 _20767_ (.A(_11326_),
    .B1(net733),
    .B2(_11424_),
    .ZN(_11431_));
 NOR2_X2 _20768_ (.A1(net162),
    .A2(_11382_),
    .ZN(_11432_));
 OAI21_X1 _20769_ (.A(_11181_),
    .B1(_11303_),
    .B2(net562),
    .ZN(_11433_));
 NOR2_X1 _20770_ (.A1(_11432_),
    .A2(_11433_),
    .ZN(_11434_));
 OR2_X1 _20771_ (.A1(_11431_),
    .A2(_11434_),
    .ZN(_11435_));
 AOI221_X2 _20772_ (.A(_11423_),
    .B1(_11430_),
    .B2(_11319_),
    .C1(_11435_),
    .C2(_11404_),
    .ZN(_11436_));
 CLKBUF_X3 _20773_ (.A(_11336_),
    .Z(_11437_));
 OAI21_X4 _20774_ (.A(_11402_),
    .B1(_11231_),
    .B2(_11235_),
    .ZN(_11438_));
 NAND3_X4 _20775_ (.A1(_11155_),
    .A2(_11278_),
    .A3(_11274_),
    .ZN(_11439_));
 OAI21_X1 _20776_ (.A(_11438_),
    .B1(_11439_),
    .B2(net511),
    .ZN(_11440_));
 AOI221_X1 _20777_ (.A(_11289_),
    .B1(_11354_),
    .B2(_11179_),
    .C1(_11440_),
    .C2(_11181_),
    .ZN(_11441_));
 INV_X2 _20778_ (.A(_14892_),
    .ZN(_11442_));
 NAND2_X1 _20779_ (.A1(_11442_),
    .A2(_11239_),
    .ZN(_11443_));
 AOI21_X2 _20780_ (.A(_11180_),
    .B1(_11285_),
    .B2(net649),
    .ZN(_11444_));
 AOI221_X1 _20781_ (.A(_11269_),
    .B1(_11352_),
    .B2(_11382_),
    .C1(_11443_),
    .C2(_11444_),
    .ZN(_11445_));
 OR3_X1 _20782_ (.A1(_11437_),
    .A2(_11441_),
    .A3(_11445_),
    .ZN(_11446_));
 NAND3_X4 _20783_ (.A1(_14906_),
    .A2(_11346_),
    .A3(_11347_),
    .ZN(_11447_));
 NAND2_X1 _20784_ (.A1(_11438_),
    .A2(_11447_),
    .ZN(_11448_));
 INV_X1 _20785_ (.A(_11129_),
    .ZN(_11449_));
 NAND2_X1 _20786_ (.A1(_06619_),
    .A2(_11207_),
    .ZN(_11450_));
 NAND2_X1 _20787_ (.A1(_11111_),
    .A2(_11207_),
    .ZN(_11451_));
 MUX2_X1 _20788_ (.A(_11450_),
    .B(_11451_),
    .S(_11125_),
    .Z(_11452_));
 AOI21_X4 _20789_ (.A(_11179_),
    .B1(_11449_),
    .B2(_11452_),
    .ZN(_11453_));
 NAND2_X1 _20790_ (.A1(_11286_),
    .A2(_11453_),
    .ZN(_11454_));
 NOR3_X4 _20791_ (.A1(_14894_),
    .A2(_11230_),
    .A3(_11234_),
    .ZN(_11455_));
 NOR3_X1 _20792_ (.A1(_11181_),
    .A2(_11289_),
    .A3(_11455_),
    .ZN(_11456_));
 AOI221_X1 _20793_ (.A(_11390_),
    .B1(_11409_),
    .B2(_11448_),
    .C1(_11454_),
    .C2(_11456_),
    .ZN(_11457_));
 AOI21_X1 _20794_ (.A(_11182_),
    .B1(_11439_),
    .B2(_11366_),
    .ZN(_11458_));
 AOI21_X1 _20795_ (.A(_11455_),
    .B1(_11374_),
    .B2(_11322_),
    .ZN(_11459_));
 AOI21_X1 _20796_ (.A(_11458_),
    .B1(_11459_),
    .B2(_14908_),
    .ZN(_11460_));
 OAI21_X1 _20797_ (.A(_11457_),
    .B1(_11460_),
    .B2(_11318_),
    .ZN(_11461_));
 NAND3_X1 _20798_ (.A1(_11358_),
    .A2(_11446_),
    .A3(_11461_),
    .ZN(_11462_));
 AOI221_X2 _20799_ (.A(_11285_),
    .B1(_11279_),
    .B2(_11131_),
    .C1(_11331_),
    .C2(_11341_),
    .ZN(_11463_));
 NOR3_X1 _20800_ (.A1(_14916_),
    .A2(_11391_),
    .A3(_11413_),
    .ZN(_11464_));
 NOR3_X1 _20801_ (.A1(_11437_),
    .A2(_11463_),
    .A3(_11464_),
    .ZN(_11465_));
 NOR2_X1 _20802_ (.A1(_11358_),
    .A2(_11465_),
    .ZN(_11466_));
 OR2_X4 _20803_ (.A1(net575),
    .A2(_11239_),
    .ZN(_11467_));
 NAND3_X1 _20804_ (.A1(_11409_),
    .A2(_11439_),
    .A3(_11467_),
    .ZN(_11468_));
 XNOR2_X1 _20805_ (.A(_11131_),
    .B(_11239_),
    .ZN(_11469_));
 OR3_X1 _20806_ (.A1(_11182_),
    .A2(_11391_),
    .A3(_11469_),
    .ZN(_11470_));
 NOR2_X2 _20807_ (.A1(_11155_),
    .A2(_11176_),
    .ZN(_11471_));
 OR4_X1 _20808_ (.A1(net162),
    .A2(_11303_),
    .A3(_11408_),
    .A4(_11471_),
    .ZN(_11472_));
 NOR2_X1 _20809_ (.A1(_11442_),
    .A2(_11326_),
    .ZN(_11473_));
 OAI21_X1 _20810_ (.A(_11304_),
    .B1(_11471_),
    .B2(_11473_),
    .ZN(_11474_));
 NAND3_X1 _20811_ (.A1(_11290_),
    .A2(_11472_),
    .A3(_11474_),
    .ZN(_11475_));
 NAND4_X1 _20812_ (.A1(_11437_),
    .A2(_11468_),
    .A3(_11470_),
    .A4(_11475_),
    .ZN(_11476_));
 AOI21_X1 _20813_ (.A(_11194_),
    .B1(_11466_),
    .B2(_11476_),
    .ZN(_11477_));
 NOR2_X2 _20814_ (.A1(_11388_),
    .A2(_11210_),
    .ZN(_11478_));
 AOI21_X1 _20815_ (.A(_11317_),
    .B1(_11307_),
    .B2(_11134_),
    .ZN(_11479_));
 INV_X1 _20816_ (.A(_14906_),
    .ZN(_11480_));
 NOR2_X2 _20817_ (.A1(_11480_),
    .A2(_11303_),
    .ZN(_11481_));
 OAI221_X1 _20818_ (.A(_11479_),
    .B1(_11481_),
    .B2(_11182_),
    .C1(_11134_),
    .C2(_11236_),
    .ZN(_11482_));
 NAND2_X1 _20819_ (.A1(_11237_),
    .A2(_11351_),
    .ZN(_11483_));
 OAI21_X1 _20820_ (.A(_11438_),
    .B1(_11373_),
    .B2(_11322_),
    .ZN(_11484_));
 OAI221_X1 _20821_ (.A(_11317_),
    .B1(_11307_),
    .B2(_11483_),
    .C1(_11484_),
    .C2(_11332_),
    .ZN(_11485_));
 AND2_X1 _20822_ (.A1(_11482_),
    .A2(_11485_),
    .ZN(_11486_));
 OAI222_X2 _20823_ (.A1(net161),
    .A2(_11428_),
    .B1(_11401_),
    .B2(_14899_),
    .C1(_11323_),
    .C2(net651),
    .ZN(_11487_));
 AOI21_X1 _20824_ (.A(_11237_),
    .B1(_11424_),
    .B2(_11438_),
    .ZN(_11488_));
 NOR2_X2 _20825_ (.A1(_11303_),
    .A2(_11453_),
    .ZN(_11489_));
 AOI21_X1 _20826_ (.A(_11488_),
    .B1(_11489_),
    .B2(_11332_),
    .ZN(_11490_));
 MUX2_X1 _20827_ (.A(_11487_),
    .B(_11490_),
    .S(_11290_),
    .Z(_11491_));
 MUX2_X1 _20828_ (.A(_11486_),
    .B(_11491_),
    .S(_11329_),
    .Z(_11492_));
 AOI221_X2 _20829_ (.A(_11436_),
    .B1(_11462_),
    .B2(_11477_),
    .C1(_11478_),
    .C2(_11492_),
    .ZN(_00057_));
 NAND2_X1 _20830_ (.A1(_14911_),
    .A2(_11297_),
    .ZN(_11493_));
 NAND2_X1 _20831_ (.A1(_11155_),
    .A2(_11176_),
    .ZN(_11494_));
 NAND3_X1 _20832_ (.A1(_14896_),
    .A2(_11319_),
    .A3(_11494_),
    .ZN(_11495_));
 NAND3_X1 _20833_ (.A1(_11287_),
    .A2(_11493_),
    .A3(_11495_),
    .ZN(_11496_));
 OAI211_X2 _20834_ (.A(_11179_),
    .B(_11331_),
    .C1(_11126_),
    .C2(_11129_),
    .ZN(_11497_));
 MUX2_X1 _20835_ (.A(_14920_),
    .B(_11497_),
    .S(_11390_),
    .Z(_11498_));
 NAND2_X1 _20836_ (.A1(_11414_),
    .A2(_11498_),
    .ZN(_11499_));
 NAND4_X1 _20837_ (.A1(_11318_),
    .A2(_11419_),
    .A3(_11496_),
    .A4(_11499_),
    .ZN(_11500_));
 NAND2_X1 _20838_ (.A1(_11292_),
    .A2(_11419_),
    .ZN(_11501_));
 NOR2_X1 _20839_ (.A1(_11286_),
    .A2(_11453_),
    .ZN(_11502_));
 NOR2_X1 _20840_ (.A1(_11283_),
    .A2(_11214_),
    .ZN(_11503_));
 OAI21_X1 _20841_ (.A(_11406_),
    .B1(_11413_),
    .B2(_11503_),
    .ZN(_11504_));
 OAI21_X1 _20842_ (.A(_11332_),
    .B1(_11374_),
    .B2(_11341_),
    .ZN(_11505_));
 OAI221_X1 _20843_ (.A(_11437_),
    .B1(_11502_),
    .B2(_11504_),
    .C1(_11505_),
    .C2(_11489_),
    .ZN(_11506_));
 OAI21_X2 _20844_ (.A(_11366_),
    .B1(_11286_),
    .B2(_11322_),
    .ZN(_11507_));
 AOI22_X1 _20845_ (.A1(_11214_),
    .A2(_11378_),
    .B1(_11507_),
    .B2(_11327_),
    .ZN(_11508_));
 OAI21_X1 _20846_ (.A(_11506_),
    .B1(_11508_),
    .B2(_11405_),
    .ZN(_11509_));
 OAI21_X1 _20847_ (.A(_11500_),
    .B1(_11501_),
    .B2(_11509_),
    .ZN(_11510_));
 OAI21_X4 _20848_ (.A(_11367_),
    .B1(_11231_),
    .B2(_11235_),
    .ZN(_11511_));
 AOI21_X1 _20849_ (.A(_11332_),
    .B1(_11439_),
    .B2(_11511_),
    .ZN(_11512_));
 NOR3_X4 _20850_ (.A1(_14906_),
    .A2(_11231_),
    .A3(_11235_),
    .ZN(_11513_));
 NOR2_X2 _20851_ (.A1(_11326_),
    .A2(_11513_),
    .ZN(_11514_));
 NAND2_X1 _20852_ (.A1(_11134_),
    .A2(_11374_),
    .ZN(_11515_));
 AOI21_X1 _20853_ (.A(_11512_),
    .B1(_11514_),
    .B2(_11515_),
    .ZN(_11516_));
 AOI21_X1 _20854_ (.A(_11316_),
    .B1(_11384_),
    .B2(_11516_),
    .ZN(_11517_));
 NAND3_X1 _20855_ (.A1(_11327_),
    .A2(_11323_),
    .A3(_11369_),
    .ZN(_11518_));
 NAND3_X1 _20856_ (.A1(_11178_),
    .A2(_11351_),
    .A3(_11447_),
    .ZN(_11519_));
 NAND2_X1 _20857_ (.A1(_11518_),
    .A2(_11519_),
    .ZN(_11520_));
 NAND3_X1 _20858_ (.A1(_11405_),
    .A2(_11318_),
    .A3(_11520_),
    .ZN(_11521_));
 NAND3_X1 _20859_ (.A1(_11332_),
    .A2(_11369_),
    .A3(_11438_),
    .ZN(_11522_));
 NAND3_X1 _20860_ (.A1(_11327_),
    .A2(_11439_),
    .A3(_11366_),
    .ZN(_11523_));
 NAND3_X1 _20861_ (.A1(_11291_),
    .A2(_11522_),
    .A3(_11523_),
    .ZN(_11524_));
 AND2_X1 _20862_ (.A1(_11214_),
    .A2(_11237_),
    .ZN(_11525_));
 OAI21_X1 _20863_ (.A(_11369_),
    .B1(_11413_),
    .B2(_11420_),
    .ZN(_11526_));
 AOI21_X1 _20864_ (.A(_11525_),
    .B1(_11526_),
    .B2(_11327_),
    .ZN(_11527_));
 OAI21_X1 _20865_ (.A(_11524_),
    .B1(_11527_),
    .B2(_11291_),
    .ZN(_11528_));
 OAI211_X2 _20866_ (.A(_11517_),
    .B(_11521_),
    .C1(_11405_),
    .C2(_11528_),
    .ZN(_11529_));
 AOI21_X2 _20867_ (.A(_11176_),
    .B1(_11239_),
    .B2(net509),
    .ZN(_11530_));
 NAND2_X1 _20868_ (.A1(net649),
    .A2(_11360_),
    .ZN(_11531_));
 AOI221_X2 _20869_ (.A(_11289_),
    .B1(_11467_),
    .B2(_11345_),
    .C1(_11530_),
    .C2(_11531_),
    .ZN(_11532_));
 OAI33_X1 _20870_ (.A1(_14906_),
    .A2(_11331_),
    .A3(_11303_),
    .B1(_11307_),
    .B2(_11282_),
    .B3(_11361_),
    .ZN(_11533_));
 AOI21_X2 _20871_ (.A(_11532_),
    .B1(_11533_),
    .B2(_11391_),
    .ZN(_11534_));
 NOR2_X1 _20872_ (.A1(_11357_),
    .A2(_11336_),
    .ZN(_11535_));
 AOI21_X1 _20873_ (.A(_11215_),
    .B1(_11323_),
    .B2(_11447_),
    .ZN(_11536_));
 AND2_X1 _20874_ (.A1(_14897_),
    .A2(_11400_),
    .ZN(_11537_));
 NOR4_X1 _20875_ (.A1(_11391_),
    .A2(_11240_),
    .A3(_11536_),
    .A4(_11537_),
    .ZN(_11538_));
 NAND2_X2 _20876_ (.A1(_11210_),
    .A2(_11336_),
    .ZN(_11539_));
 NOR2_X1 _20877_ (.A1(_11538_),
    .A2(_11539_),
    .ZN(_11540_));
 OR2_X2 _20878_ (.A1(_11344_),
    .A2(_11331_),
    .ZN(_11541_));
 OAI21_X1 _20879_ (.A(_11177_),
    .B1(_11413_),
    .B2(_11283_),
    .ZN(_11542_));
 NOR2_X2 _20880_ (.A1(net162),
    .A2(_11373_),
    .ZN(_11543_));
 OAI221_X2 _20881_ (.A(_11290_),
    .B1(_11541_),
    .B2(_11361_),
    .C1(_11542_),
    .C2(_11543_),
    .ZN(_11544_));
 AOI221_X2 _20882_ (.A(_11194_),
    .B1(_11535_),
    .B2(_11534_),
    .C1(_11540_),
    .C2(_11544_),
    .ZN(_11545_));
 OAI211_X2 _20883_ (.A(_11406_),
    .B(_11343_),
    .C1(_11286_),
    .C2(_11420_),
    .ZN(_11546_));
 OAI21_X1 _20884_ (.A(_11546_),
    .B1(_11507_),
    .B2(_11182_),
    .ZN(_11547_));
 NAND2_X2 _20885_ (.A1(_11155_),
    .A2(_11215_),
    .ZN(_11548_));
 NAND3_X1 _20886_ (.A1(_11420_),
    .A2(_11286_),
    .A3(_11548_),
    .ZN(_11549_));
 NAND2_X1 _20887_ (.A1(_11133_),
    .A2(_11326_),
    .ZN(_11550_));
 MUX2_X1 _20888_ (.A(_11215_),
    .B(_11373_),
    .S(_11131_),
    .Z(_11551_));
 OAI221_X1 _20889_ (.A(_11549_),
    .B1(_11550_),
    .B2(_11348_),
    .C1(net161),
    .C2(_11551_),
    .ZN(_11552_));
 MUX2_X1 _20890_ (.A(_11547_),
    .B(_11552_),
    .S(_11290_),
    .Z(_11553_));
 NOR2_X2 _20891_ (.A1(_11312_),
    .A2(_11215_),
    .ZN(_11554_));
 NOR2_X1 _20892_ (.A1(_11308_),
    .A2(_11155_),
    .ZN(_11555_));
 AOI221_X2 _20893_ (.A(_11554_),
    .B1(_11347_),
    .B2(_11346_),
    .C1(_11406_),
    .C2(_11555_),
    .ZN(_11556_));
 AOI21_X1 _20894_ (.A(_11317_),
    .B1(_11304_),
    .B2(_14913_),
    .ZN(_11557_));
 INV_X1 _20895_ (.A(_11557_),
    .ZN(_11558_));
 AOI221_X2 _20896_ (.A(_11411_),
    .B1(_11347_),
    .B2(_11346_),
    .C1(net651),
    .C2(_11326_),
    .ZN(_11559_));
 OAI21_X1 _20897_ (.A(_11299_),
    .B1(_11287_),
    .B2(_14916_),
    .ZN(_11560_));
 OAI22_X1 _20898_ (.A1(_11556_),
    .A2(_11558_),
    .B1(_11559_),
    .B2(_11560_),
    .ZN(_11561_));
 MUX2_X1 _20899_ (.A(_11553_),
    .B(_11561_),
    .S(_11329_),
    .Z(_11562_));
 AOI221_X2 _20900_ (.A(_11510_),
    .B1(_11545_),
    .B2(_11529_),
    .C1(_11562_),
    .C2(_11478_),
    .ZN(_00058_));
 INV_X1 _20901_ (.A(_11419_),
    .ZN(_11563_));
 NAND3_X1 _20902_ (.A1(_11327_),
    .A2(_11319_),
    .A3(_11287_),
    .ZN(_11564_));
 NOR3_X4 _20903_ (.A1(_11180_),
    .A2(_11295_),
    .A3(_11257_),
    .ZN(_11565_));
 NAND2_X1 _20904_ (.A1(_14896_),
    .A2(_11565_),
    .ZN(_11566_));
 OAI221_X1 _20905_ (.A(_11564_),
    .B1(_11565_),
    .B2(net733),
    .C1(_11330_),
    .C2(_11566_),
    .ZN(_11567_));
 NAND3_X1 _20906_ (.A1(net196),
    .A2(_11414_),
    .A3(_11548_),
    .ZN(_11568_));
 AOI21_X1 _20907_ (.A(_11319_),
    .B1(_11408_),
    .B2(_14896_),
    .ZN(_11569_));
 AOI21_X1 _20908_ (.A(_11279_),
    .B1(_11354_),
    .B2(_14896_),
    .ZN(_11570_));
 AOI22_X1 _20909_ (.A1(_11568_),
    .A2(_11569_),
    .B1(_11570_),
    .B2(_11437_),
    .ZN(_11571_));
 OR3_X1 _20910_ (.A1(_11292_),
    .A2(_11567_),
    .A3(_11571_),
    .ZN(_11572_));
 NAND2_X1 _20911_ (.A1(_11406_),
    .A2(_11336_),
    .ZN(_11573_));
 NAND2_X1 _20912_ (.A1(_11341_),
    .A2(_11304_),
    .ZN(_11574_));
 AOI21_X1 _20913_ (.A(_11573_),
    .B1(_11574_),
    .B2(_11397_),
    .ZN(_11575_));
 AOI21_X4 _20914_ (.A(_11215_),
    .B1(_11254_),
    .B2(_11258_),
    .ZN(_11576_));
 NOR2_X1 _20915_ (.A1(net734),
    .A2(_11413_),
    .ZN(_11577_));
 NOR2_X1 _20916_ (.A1(_11307_),
    .A2(_11577_),
    .ZN(_11578_));
 OAI22_X2 _20917_ (.A1(_11541_),
    .A2(_11481_),
    .B1(_11483_),
    .B2(_11543_),
    .ZN(_11579_));
 AOI221_X1 _20918_ (.A(_11575_),
    .B1(_11576_),
    .B2(_11578_),
    .C1(_11579_),
    .C2(_11329_),
    .ZN(_11580_));
 OAI21_X1 _20919_ (.A(_11572_),
    .B1(_11580_),
    .B2(_11300_),
    .ZN(_11581_));
 AOI22_X1 _20920_ (.A1(_11283_),
    .A2(_11287_),
    .B1(_11344_),
    .B2(_11290_),
    .ZN(_11582_));
 OR2_X1 _20921_ (.A1(_14915_),
    .A2(_11582_),
    .ZN(_11583_));
 NAND4_X1 _20922_ (.A1(_14915_),
    .A2(_11300_),
    .A3(net733),
    .A4(_11574_),
    .ZN(_11584_));
 BUF_X16 _20923_ (.A(_11376_),
    .Z(_14891_));
 NAND3_X1 _20924_ (.A1(net197),
    .A2(_11300_),
    .A3(_11400_),
    .ZN(_11585_));
 NAND4_X1 _20925_ (.A1(_11405_),
    .A2(_11583_),
    .A3(_11584_),
    .A4(_11585_),
    .ZN(_11586_));
 AOI22_X2 _20926_ (.A1(_11368_),
    .A2(_11401_),
    .B1(_11279_),
    .B2(_11304_),
    .ZN(_11587_));
 OAI21_X1 _20927_ (.A(_11333_),
    .B1(_11307_),
    .B2(_11481_),
    .ZN(_11588_));
 NAND2_X1 _20928_ (.A1(_11390_),
    .A2(_11317_),
    .ZN(_11589_));
 NAND2_X1 _20929_ (.A1(_11374_),
    .A2(_11503_),
    .ZN(_11590_));
 AOI21_X1 _20930_ (.A(_11589_),
    .B1(_11393_),
    .B2(_11590_),
    .ZN(_11591_));
 AOI221_X2 _20931_ (.A(_11194_),
    .B1(_11270_),
    .B2(_11587_),
    .C1(_11588_),
    .C2(_11591_),
    .ZN(_11592_));
 AOI21_X1 _20932_ (.A(_11358_),
    .B1(_11586_),
    .B2(_11592_),
    .ZN(_11593_));
 AOI221_X2 _20933_ (.A(_11259_),
    .B1(_11310_),
    .B2(_11442_),
    .C1(_11353_),
    .C2(net649),
    .ZN(_11594_));
 OAI21_X1 _20934_ (.A(_11594_),
    .B1(_11530_),
    .B2(_14890_),
    .ZN(_11595_));
 NAND3_X4 _20935_ (.A1(_11347_),
    .A2(_11346_),
    .A3(net10),
    .ZN(_11596_));
 AND2_X1 _20936_ (.A1(_11511_),
    .A2(_11596_),
    .ZN(_11597_));
 NAND3_X1 _20937_ (.A1(_11182_),
    .A2(_11319_),
    .A3(_11597_),
    .ZN(_11598_));
 NAND3_X1 _20938_ (.A1(_11375_),
    .A2(_11447_),
    .A3(_11576_),
    .ZN(_11599_));
 NOR2_X2 _20939_ (.A1(_11194_),
    .A2(_11317_),
    .ZN(_11600_));
 AND4_X1 _20940_ (.A1(_11595_),
    .A2(_11598_),
    .A3(_11599_),
    .A4(_11600_),
    .ZN(_11601_));
 NOR2_X1 _20941_ (.A1(net562),
    .A2(_11181_),
    .ZN(_11602_));
 OAI21_X1 _20942_ (.A(_11336_),
    .B1(_11413_),
    .B2(_11602_),
    .ZN(_11603_));
 NOR2_X1 _20943_ (.A1(_11413_),
    .A2(_11565_),
    .ZN(_11604_));
 AOI21_X1 _20944_ (.A(_11307_),
    .B1(_11336_),
    .B2(_11420_),
    .ZN(_11605_));
 OAI221_X1 _20945_ (.A(_11603_),
    .B1(_11604_),
    .B2(_11335_),
    .C1(_11178_),
    .C2(_11605_),
    .ZN(_11606_));
 NOR2_X1 _20946_ (.A1(_11390_),
    .A2(_11286_),
    .ZN(_11607_));
 NAND2_X1 _20947_ (.A1(_11368_),
    .A2(_11237_),
    .ZN(_11608_));
 OAI21_X1 _20948_ (.A(_11608_),
    .B1(_11177_),
    .B2(_11312_),
    .ZN(_11609_));
 AOI21_X1 _20949_ (.A(_11290_),
    .B1(_11607_),
    .B2(_11609_),
    .ZN(_11610_));
 AOI21_X1 _20950_ (.A(_11388_),
    .B1(_11606_),
    .B2(_11610_),
    .ZN(_11611_));
 AOI221_X1 _20951_ (.A(_11259_),
    .B1(_11310_),
    .B2(_11341_),
    .C1(_11354_),
    .C2(_11402_),
    .ZN(_11612_));
 AOI22_X1 _20952_ (.A1(_14899_),
    .A2(_11400_),
    .B1(_11272_),
    .B2(_11286_),
    .ZN(_11613_));
 OAI21_X1 _20953_ (.A(_11612_),
    .B1(_11613_),
    .B2(net196),
    .ZN(_11614_));
 NOR2_X1 _20954_ (.A1(_11342_),
    .A2(_11180_),
    .ZN(_11615_));
 AOI221_X1 _20955_ (.A(_11296_),
    .B1(_11239_),
    .B2(_11615_),
    .C1(_11361_),
    .C2(_11308_),
    .ZN(_11616_));
 OAI21_X1 _20956_ (.A(_11616_),
    .B1(_11541_),
    .B2(_11361_),
    .ZN(_11617_));
 NAND3_X1 _20957_ (.A1(_11617_),
    .A2(_11614_),
    .A3(_11291_),
    .ZN(_11618_));
 OAI221_X1 _20958_ (.A(_11304_),
    .B1(_11257_),
    .B2(_11295_),
    .C1(_11480_),
    .C2(_11406_),
    .ZN(_11619_));
 OAI21_X1 _20959_ (.A(_11299_),
    .B1(_11279_),
    .B2(_11619_),
    .ZN(_11620_));
 INV_X1 _20960_ (.A(_11367_),
    .ZN(_11621_));
 NAND2_X1 _20961_ (.A1(_11207_),
    .A2(_11621_),
    .ZN(_11622_));
 NOR3_X1 _20962_ (.A1(_11156_),
    .A2(_11167_),
    .A3(_11160_),
    .ZN(_11623_));
 XNOR2_X1 _20963_ (.A(_11167_),
    .B(_11162_),
    .ZN(_11624_));
 AOI21_X1 _20964_ (.A(_11623_),
    .B1(_11624_),
    .B2(_11156_),
    .ZN(_11625_));
 OAI22_X1 _20965_ (.A1(_11231_),
    .A2(_11235_),
    .B1(_11622_),
    .B2(_11625_),
    .ZN(_11626_));
 OR2_X4 _20966_ (.A1(_14897_),
    .A2(_14894_),
    .ZN(_11627_));
 XNOR2_X1 _20967_ (.A(_06635_),
    .B(_00451_),
    .ZN(_11628_));
 MUX2_X1 _20968_ (.A(_11368_),
    .B(_11627_),
    .S(_11628_),
    .Z(_11629_));
 NAND2_X1 _20969_ (.A1(_09136_),
    .A2(_11629_),
    .ZN(_11630_));
 NOR3_X1 _20970_ (.A1(_11156_),
    .A2(_11367_),
    .A3(_11162_),
    .ZN(_11631_));
 AOI21_X1 _20971_ (.A(_09136_),
    .B1(_11167_),
    .B2(_11631_),
    .ZN(_11632_));
 XNOR2_X1 _20972_ (.A(_11156_),
    .B(_11624_),
    .ZN(_11633_));
 OAI21_X1 _20973_ (.A(_11632_),
    .B1(_11633_),
    .B2(_11627_),
    .ZN(_11634_));
 AOI21_X1 _20974_ (.A(_11626_),
    .B1(_11630_),
    .B2(_11634_),
    .ZN(_11635_));
 NOR3_X1 _20975_ (.A1(_11635_),
    .A2(_11463_),
    .A3(_11319_),
    .ZN(_11636_));
 OAI21_X1 _20976_ (.A(_11358_),
    .B1(_11636_),
    .B2(_11620_),
    .ZN(_11637_));
 AOI221_X2 _20977_ (.A(_11601_),
    .B1(_11611_),
    .B2(_11618_),
    .C1(_11637_),
    .C2(_11388_),
    .ZN(_11638_));
 OAI22_X1 _20978_ (.A1(_11563_),
    .A2(_11581_),
    .B1(_11638_),
    .B2(_11593_),
    .ZN(_00059_));
 NOR2_X2 _20979_ (.A1(_11194_),
    .A2(_11357_),
    .ZN(_11639_));
 NOR2_X1 _20980_ (.A1(_11402_),
    .A2(_11215_),
    .ZN(_11640_));
 MUX2_X1 _20981_ (.A(_14904_),
    .B(_11640_),
    .S(_11373_),
    .Z(_11641_));
 OAI21_X1 _20982_ (.A(_11639_),
    .B1(_11641_),
    .B2(_11392_),
    .ZN(_11642_));
 AOI21_X1 _20983_ (.A(_11432_),
    .B1(_11511_),
    .B2(_11332_),
    .ZN(_11643_));
 NAND2_X1 _20984_ (.A1(_11336_),
    .A2(_11391_),
    .ZN(_11644_));
 AOI21_X1 _20985_ (.A(_11644_),
    .B1(_11310_),
    .B2(net196),
    .ZN(_11645_));
 AOI21_X1 _20986_ (.A(_11360_),
    .B1(_11239_),
    .B2(net509),
    .ZN(_11646_));
 NAND2_X1 _20987_ (.A1(_11176_),
    .A2(_11285_),
    .ZN(_11647_));
 OAI221_X1 _20988_ (.A(_11396_),
    .B1(_11646_),
    .B2(_11331_),
    .C1(_11647_),
    .C2(_11621_),
    .ZN(_11648_));
 AOI22_X1 _20989_ (.A1(_11442_),
    .A2(_11354_),
    .B1(_11361_),
    .B2(net510),
    .ZN(_11649_));
 OAI21_X1 _20990_ (.A(_11649_),
    .B1(_11325_),
    .B2(_11237_),
    .ZN(_11650_));
 MUX2_X1 _20991_ (.A(_11648_),
    .B(_11650_),
    .S(_11390_),
    .Z(_11651_));
 AOI221_X2 _20992_ (.A(_11642_),
    .B1(_11643_),
    .B2(_11645_),
    .C1(_11651_),
    .C2(_11299_),
    .ZN(_11652_));
 AOI21_X2 _20993_ (.A(_11554_),
    .B1(_11182_),
    .B2(_11214_),
    .ZN(_11653_));
 AOI221_X2 _20994_ (.A(_11317_),
    .B1(_11455_),
    .B2(_11576_),
    .C1(_11653_),
    .C2(_11281_),
    .ZN(_11654_));
 NAND2_X1 _20995_ (.A1(_14890_),
    .A2(_11565_),
    .ZN(_11655_));
 OAI21_X1 _20996_ (.A(_11453_),
    .B1(_11337_),
    .B2(_11576_),
    .ZN(_11656_));
 AND2_X1 _20997_ (.A1(_11655_),
    .A2(_11656_),
    .ZN(_11657_));
 OAI21_X1 _20998_ (.A(_11654_),
    .B1(_11657_),
    .B2(_11330_),
    .ZN(_11658_));
 AOI221_X1 _20999_ (.A(_11259_),
    .B1(_11354_),
    .B2(_11480_),
    .C1(_11382_),
    .C2(_11326_),
    .ZN(_11659_));
 AOI221_X1 _21000_ (.A(_11296_),
    .B1(_11352_),
    .B2(_11443_),
    .C1(_11469_),
    .C2(_11237_),
    .ZN(_11660_));
 OAI21_X1 _21001_ (.A(_11318_),
    .B1(_11659_),
    .B2(_11660_),
    .ZN(_11661_));
 AND2_X1 _21002_ (.A1(_11211_),
    .A2(_11661_),
    .ZN(_11662_));
 NAND2_X1 _21003_ (.A1(_14892_),
    .A2(_11239_),
    .ZN(_11663_));
 AOI221_X2 _21004_ (.A(_11259_),
    .B1(_11663_),
    .B2(_11444_),
    .C1(_11326_),
    .C2(_11155_),
    .ZN(_11664_));
 AOI21_X1 _21005_ (.A(_11455_),
    .B1(_11511_),
    .B2(_11177_),
    .ZN(_11665_));
 NOR2_X1 _21006_ (.A1(_11297_),
    .A2(_11665_),
    .ZN(_11666_));
 NOR4_X1 _21007_ (.A1(_11316_),
    .A2(_11318_),
    .A3(_11664_),
    .A4(_11666_),
    .ZN(_11667_));
 NAND3_X1 _21008_ (.A1(_11134_),
    .A2(_11406_),
    .A3(_11390_),
    .ZN(_11668_));
 NAND2_X1 _21009_ (.A1(_11322_),
    .A2(_11576_),
    .ZN(_11669_));
 AOI21_X1 _21010_ (.A(_11304_),
    .B1(_11668_),
    .B2(_11669_),
    .ZN(_11670_));
 OAI21_X1 _21011_ (.A(net651),
    .B1(_14899_),
    .B2(_11565_),
    .ZN(_11671_));
 AOI21_X1 _21012_ (.A(_11374_),
    .B1(_11548_),
    .B2(_11671_),
    .ZN(_11672_));
 AOI21_X1 _21013_ (.A(_11134_),
    .B1(_11362_),
    .B2(_11573_),
    .ZN(_11673_));
 NOR4_X2 _21014_ (.A1(_11359_),
    .A2(_11670_),
    .A3(_11672_),
    .A4(_11673_),
    .ZN(_11674_));
 NOR2_X1 _21015_ (.A1(_11621_),
    .A2(_11177_),
    .ZN(_11675_));
 NOR3_X1 _21016_ (.A1(_11299_),
    .A2(_11431_),
    .A3(_11675_),
    .ZN(_11676_));
 NOR2_X1 _21017_ (.A1(_11176_),
    .A2(_11363_),
    .ZN(_11677_));
 AOI21_X2 _21018_ (.A(_11513_),
    .B1(_11285_),
    .B2(_11308_),
    .ZN(_11678_));
 AOI221_X2 _21019_ (.A(_11289_),
    .B1(_11531_),
    .B2(_11677_),
    .C1(_11678_),
    .C2(_11237_),
    .ZN(_11679_));
 NOR3_X1 _21020_ (.A1(_11539_),
    .A2(_11676_),
    .A3(_11679_),
    .ZN(_11680_));
 NOR4_X1 _21021_ (.A1(_11680_),
    .A2(_11667_),
    .A3(_11674_),
    .A4(_11388_),
    .ZN(_11681_));
 NAND2_X1 _21022_ (.A1(_14908_),
    .A2(_11397_),
    .ZN(_11682_));
 OR2_X1 _21023_ (.A1(_11240_),
    .A2(_11363_),
    .ZN(_11683_));
 OAI221_X2 _21024_ (.A(_11300_),
    .B1(_11432_),
    .B2(_11682_),
    .C1(_11683_),
    .C2(_14908_),
    .ZN(_11684_));
 NOR2_X1 _21025_ (.A1(_11308_),
    .A2(_11375_),
    .ZN(_11685_));
 OR2_X1 _21026_ (.A1(_11178_),
    .A2(_11513_),
    .ZN(_11686_));
 OAI221_X1 _21027_ (.A(_11291_),
    .B1(_11685_),
    .B2(_11686_),
    .C1(_11597_),
    .C2(_14908_),
    .ZN(_11687_));
 NAND3_X1 _21028_ (.A1(_11535_),
    .A2(_11684_),
    .A3(_11687_),
    .ZN(_11688_));
 AOI221_X1 _21029_ (.A(_11652_),
    .B1(_11658_),
    .B2(_11662_),
    .C1(_11681_),
    .C2(_11688_),
    .ZN(_00060_));
 NOR3_X1 _21030_ (.A1(_11388_),
    .A2(_11358_),
    .A3(_11318_),
    .ZN(_11689_));
 OAI21_X1 _21031_ (.A(_14891_),
    .B1(_11329_),
    .B2(_11414_),
    .ZN(_11690_));
 AOI22_X1 _21032_ (.A1(_11341_),
    .A2(_11378_),
    .B1(_11400_),
    .B2(_14890_),
    .ZN(_11691_));
 OAI221_X1 _21033_ (.A(_11689_),
    .B1(_11690_),
    .B2(_11354_),
    .C1(_11691_),
    .C2(_11298_),
    .ZN(_11692_));
 NAND2_X1 _21034_ (.A1(_11405_),
    .A2(_11330_),
    .ZN(_11693_));
 AOI21_X1 _21035_ (.A(net197),
    .B1(_11329_),
    .B2(_11330_),
    .ZN(_11694_));
 AOI22_X1 _21036_ (.A1(net197),
    .A2(_11693_),
    .B1(_11694_),
    .B2(_11564_),
    .ZN(_11695_));
 AOI21_X1 _21037_ (.A(_11692_),
    .B1(_11695_),
    .B2(_14899_),
    .ZN(_11696_));
 NAND2_X1 _21038_ (.A1(_11291_),
    .A2(_11478_),
    .ZN(_11697_));
 AOI221_X2 _21039_ (.A(_11390_),
    .B1(_11286_),
    .B2(_11214_),
    .C1(_11354_),
    .C2(_11368_),
    .ZN(_11698_));
 AOI21_X1 _21040_ (.A(_11178_),
    .B1(_11324_),
    .B2(_11351_),
    .ZN(_11699_));
 AOI21_X1 _21041_ (.A(_11699_),
    .B1(_11309_),
    .B2(_11333_),
    .ZN(_11700_));
 AOI221_X2 _21042_ (.A(_11697_),
    .B1(_11698_),
    .B2(_11383_),
    .C1(_11298_),
    .C2(_11700_),
    .ZN(_11701_));
 NOR2_X1 _21043_ (.A1(_11696_),
    .A2(_11701_),
    .ZN(_11702_));
 OAI221_X1 _21044_ (.A(_11358_),
    .B1(_11400_),
    .B2(_14890_),
    .C1(_11361_),
    .C2(net197),
    .ZN(_11703_));
 OAI21_X1 _21045_ (.A(_11548_),
    .B1(_11238_),
    .B2(_11357_),
    .ZN(_11704_));
 NOR2_X1 _21046_ (.A1(_11357_),
    .A2(_11627_),
    .ZN(_11705_));
 AOI221_X1 _21047_ (.A(_11437_),
    .B1(_11543_),
    .B2(_11704_),
    .C1(_11705_),
    .C2(_11310_),
    .ZN(_11706_));
 AND2_X1 _21048_ (.A1(_11703_),
    .A2(_11706_),
    .ZN(_11707_));
 OAI221_X1 _21049_ (.A(_11178_),
    .B1(_11374_),
    .B2(_11368_),
    .C1(_11375_),
    .C2(_11376_),
    .ZN(_11708_));
 OAI21_X1 _21050_ (.A(net733),
    .B1(_11374_),
    .B2(_11420_),
    .ZN(_11709_));
 AOI21_X1 _21051_ (.A(_11316_),
    .B1(_11709_),
    .B2(_11327_),
    .ZN(_11710_));
 OAI22_X1 _21052_ (.A1(net562),
    .A2(_11647_),
    .B1(_11525_),
    .B2(_11287_),
    .ZN(_11711_));
 AOI221_X1 _21053_ (.A(_11329_),
    .B1(_11710_),
    .B2(_11708_),
    .C1(_11711_),
    .C2(_11316_),
    .ZN(_11712_));
 OAI21_X1 _21054_ (.A(_11600_),
    .B1(_11707_),
    .B2(_11712_),
    .ZN(_11713_));
 NAND2_X1 _21055_ (.A1(_11318_),
    .A2(_11211_),
    .ZN(_11714_));
 AOI21_X1 _21056_ (.A(_11406_),
    .B1(_11343_),
    .B2(_11447_),
    .ZN(_11715_));
 AOI21_X1 _21057_ (.A(_11715_),
    .B1(_11502_),
    .B2(_11327_),
    .ZN(_11716_));
 OAI21_X1 _21058_ (.A(_11414_),
    .B1(_11279_),
    .B2(_11525_),
    .ZN(_11717_));
 AOI221_X1 _21059_ (.A(_11714_),
    .B1(_11716_),
    .B2(_11437_),
    .C1(_11281_),
    .C2(_11717_),
    .ZN(_11718_));
 NAND2_X1 _21060_ (.A1(_11299_),
    .A2(_11639_),
    .ZN(_11719_));
 AND3_X4 _21061_ (.A1(_11596_),
    .A2(_14908_),
    .A3(_11438_),
    .ZN(_11720_));
 OAI21_X4 _21062_ (.A(_11405_),
    .B1(_11715_),
    .B2(_11720_),
    .ZN(_11721_));
 OAI221_X1 _21063_ (.A(_11298_),
    .B1(_11330_),
    .B2(_11342_),
    .C1(_11396_),
    .C2(_14915_),
    .ZN(_11722_));
 AOI21_X2 _21064_ (.A(_11719_),
    .B1(_11721_),
    .B2(_11722_),
    .ZN(_11723_));
 NAND3_X1 _21065_ (.A1(_11182_),
    .A2(_11596_),
    .A3(_11511_),
    .ZN(_11724_));
 AOI21_X1 _21066_ (.A(_11336_),
    .B1(_11378_),
    .B2(_14899_),
    .ZN(_11725_));
 AOI22_X2 _21067_ (.A1(_11134_),
    .A2(_11361_),
    .B1(_11424_),
    .B2(_11182_),
    .ZN(_11726_));
 AOI221_X2 _21068_ (.A(_11316_),
    .B1(_11724_),
    .B2(_11725_),
    .C1(_11726_),
    .C2(_11319_),
    .ZN(_11727_));
 NAND2_X1 _21069_ (.A1(_11194_),
    .A2(_11300_),
    .ZN(_11728_));
 NAND2_X2 _21070_ (.A1(_11324_),
    .A2(_11366_),
    .ZN(_11729_));
 AOI221_X2 _21071_ (.A(_11539_),
    .B1(_11729_),
    .B2(_11332_),
    .C1(_11400_),
    .C2(net196),
    .ZN(_11730_));
 NAND2_X1 _21072_ (.A1(_11210_),
    .A2(_11390_),
    .ZN(_11731_));
 AOI221_X2 _21073_ (.A(_11731_),
    .B1(_11514_),
    .B2(_11397_),
    .C1(_11402_),
    .C2(_11310_),
    .ZN(_11732_));
 NOR4_X2 _21074_ (.A1(_11727_),
    .A2(_11728_),
    .A3(_11730_),
    .A4(_11732_),
    .ZN(_11733_));
 NOR3_X2 _21075_ (.A1(_11718_),
    .A2(_11723_),
    .A3(_11733_),
    .ZN(_11734_));
 NAND3_X2 _21076_ (.A1(_11734_),
    .A2(_11713_),
    .A3(_11702_),
    .ZN(_00061_));
 NAND2_X1 _21077_ (.A1(_11376_),
    .A2(_11437_),
    .ZN(_11735_));
 AND3_X1 _21078_ (.A1(_14915_),
    .A2(_11362_),
    .A3(_11735_),
    .ZN(_11736_));
 AOI21_X1 _21079_ (.A(_11414_),
    .B1(_11297_),
    .B2(_11621_),
    .ZN(_11737_));
 NOR2_X1 _21080_ (.A1(_11437_),
    .A2(_11596_),
    .ZN(_11738_));
 NOR3_X1 _21081_ (.A1(_14915_),
    .A2(_11737_),
    .A3(_11738_),
    .ZN(_11739_));
 OAI221_X1 _21082_ (.A(_11300_),
    .B1(_11736_),
    .B2(_11739_),
    .C1(_11693_),
    .C2(_14890_),
    .ZN(_11740_));
 AOI21_X1 _21083_ (.A(_11307_),
    .B1(_11471_),
    .B2(net197),
    .ZN(_11741_));
 OAI221_X1 _21084_ (.A(_11494_),
    .B1(_11375_),
    .B2(_14896_),
    .C1(_11741_),
    .C2(net562),
    .ZN(_11742_));
 NAND3_X1 _21085_ (.A1(_11134_),
    .A2(_14890_),
    .A3(_11390_),
    .ZN(_11743_));
 OAI21_X1 _21086_ (.A(_14908_),
    .B1(_11297_),
    .B2(_11513_),
    .ZN(_11744_));
 NAND2_X1 _21087_ (.A1(_11297_),
    .A2(_11287_),
    .ZN(_11745_));
 OAI221_X1 _21088_ (.A(_11743_),
    .B1(_11744_),
    .B2(net197),
    .C1(_11548_),
    .C2(_11745_),
    .ZN(_11746_));
 AOI22_X1 _21089_ (.A1(_11384_),
    .A2(_11742_),
    .B1(_11746_),
    .B2(_11292_),
    .ZN(_11747_));
 NAND3_X1 _21090_ (.A1(_11211_),
    .A2(_11740_),
    .A3(_11747_),
    .ZN(_11748_));
 AND2_X1 _21091_ (.A1(_11382_),
    .A2(_11511_),
    .ZN(_11749_));
 AOI21_X1 _21092_ (.A(_11344_),
    .B1(_11627_),
    .B2(_11373_),
    .ZN(_11750_));
 MUX2_X1 _21093_ (.A(_11749_),
    .B(_11750_),
    .S(_11237_),
    .Z(_11751_));
 OAI21_X1 _21094_ (.A(_11511_),
    .B1(_11374_),
    .B2(_11322_),
    .ZN(_11752_));
 NAND2_X1 _21095_ (.A1(_14908_),
    .A2(_11752_),
    .ZN(_11753_));
 AOI21_X1 _21096_ (.A(_11299_),
    .B1(_11378_),
    .B2(_11283_),
    .ZN(_11754_));
 AOI221_X2 _21097_ (.A(_11297_),
    .B1(_11299_),
    .B2(_11751_),
    .C1(_11753_),
    .C2(_11754_),
    .ZN(_11755_));
 NAND2_X1 _21098_ (.A1(_11333_),
    .A2(_11369_),
    .ZN(_11756_));
 INV_X1 _21099_ (.A(_11283_),
    .ZN(_11757_));
 OAI21_X1 _21100_ (.A(_11447_),
    .B1(_11414_),
    .B2(_11757_),
    .ZN(_11758_));
 OAI221_X1 _21101_ (.A(_11404_),
    .B1(_11489_),
    .B2(_11756_),
    .C1(_11758_),
    .C2(_14915_),
    .ZN(_11759_));
 AOI221_X2 _21102_ (.A(_11453_),
    .B1(_11347_),
    .B2(_11346_),
    .C1(_11420_),
    .C2(_11326_),
    .ZN(_11760_));
 NOR3_X1 _21103_ (.A1(_14909_),
    .A2(_14918_),
    .A3(_11374_),
    .ZN(_11761_));
 OR3_X1 _21104_ (.A1(_11392_),
    .A2(_11760_),
    .A3(_11761_),
    .ZN(_11762_));
 NAND3_X1 _21105_ (.A1(_11358_),
    .A2(_11759_),
    .A3(_11762_),
    .ZN(_11763_));
 OAI21_X1 _21106_ (.A(_11194_),
    .B1(_11755_),
    .B2(_11763_),
    .ZN(_11764_));
 OR2_X1 _21107_ (.A1(_11215_),
    .A2(_11455_),
    .ZN(_11765_));
 OAI21_X4 _21108_ (.A(_11596_),
    .B1(_11303_),
    .B2(_11133_),
    .ZN(_11766_));
 OAI221_X2 _21109_ (.A(_11391_),
    .B1(_11685_),
    .B2(_11765_),
    .C1(_11766_),
    .C2(_11177_),
    .ZN(_11767_));
 OAI21_X2 _21110_ (.A(_11181_),
    .B1(_11373_),
    .B2(_11627_),
    .ZN(_11768_));
 NAND2_X1 _21111_ (.A1(_11323_),
    .A2(_11596_),
    .ZN(_11769_));
 OAI221_X1 _21112_ (.A(_11317_),
    .B1(_11685_),
    .B2(_11768_),
    .C1(_11769_),
    .C2(_11406_),
    .ZN(_11770_));
 AND2_X2 _21113_ (.A1(_11770_),
    .A2(_11767_),
    .ZN(_11771_));
 OAI21_X1 _21114_ (.A(_11286_),
    .B1(_11279_),
    .B2(_11420_),
    .ZN(_11772_));
 AND2_X1 _21115_ (.A1(_11381_),
    .A2(_11772_),
    .ZN(_11773_));
 AOI21_X1 _21116_ (.A(_11297_),
    .B1(_11318_),
    .B2(_11773_),
    .ZN(_11774_));
 OAI21_X1 _21117_ (.A(_11497_),
    .B1(_11177_),
    .B2(_11312_),
    .ZN(_11775_));
 MUX2_X1 _21118_ (.A(_14911_),
    .B(_11775_),
    .S(_11413_),
    .Z(_11776_));
 NAND2_X1 _21119_ (.A1(_11291_),
    .A2(_11776_),
    .ZN(_11777_));
 AOI221_X2 _21120_ (.A(_11358_),
    .B1(_11771_),
    .B2(_11329_),
    .C1(_11774_),
    .C2(_11777_),
    .ZN(_11778_));
 MUX2_X1 _21121_ (.A(_11214_),
    .B(_11368_),
    .S(_11259_),
    .Z(_11779_));
 AOI21_X1 _21122_ (.A(_11177_),
    .B1(_11336_),
    .B2(_11420_),
    .ZN(_11780_));
 AOI22_X2 _21123_ (.A1(_11333_),
    .A2(_11779_),
    .B1(_11780_),
    .B2(_11743_),
    .ZN(_11781_));
 AOI221_X2 _21124_ (.A(_11291_),
    .B1(_11615_),
    .B2(_11607_),
    .C1(_11781_),
    .C2(_11287_),
    .ZN(_11782_));
 NOR2_X1 _21125_ (.A1(_14910_),
    .A2(_11414_),
    .ZN(_11783_));
 OAI21_X1 _21126_ (.A(_11608_),
    .B1(_14915_),
    .B2(net197),
    .ZN(_11784_));
 AOI21_X1 _21127_ (.A(_11783_),
    .B1(_11784_),
    .B2(_11330_),
    .ZN(_11785_));
 AOI21_X1 _21128_ (.A(_11329_),
    .B1(_11310_),
    .B2(net161),
    .ZN(_11786_));
 AOI22_X1 _21129_ (.A1(_11298_),
    .A2(_11785_),
    .B1(_11786_),
    .B2(_11588_),
    .ZN(_11787_));
 AOI21_X1 _21130_ (.A(_11782_),
    .B1(_11787_),
    .B2(_11292_),
    .ZN(_11788_));
 OAI221_X1 _21131_ (.A(_11748_),
    .B1(_11778_),
    .B2(_11764_),
    .C1(_11389_),
    .C2(_11788_),
    .ZN(_00062_));
 NAND2_X1 _21132_ (.A1(_11405_),
    .A2(_11478_),
    .ZN(_11789_));
 NAND3_X1 _21133_ (.A1(_11333_),
    .A2(_11382_),
    .A3(_11511_),
    .ZN(_11790_));
 AOI21_X1 _21134_ (.A(_11301_),
    .B1(_11504_),
    .B2(_11790_),
    .ZN(_11791_));
 NOR2_X1 _21135_ (.A1(_11300_),
    .A2(_11791_),
    .ZN(_11792_));
 NOR3_X1 _21136_ (.A1(_11292_),
    .A2(_11363_),
    .A3(_11760_),
    .ZN(_11793_));
 AOI22_X1 _21137_ (.A1(_11480_),
    .A2(_11310_),
    .B1(_11354_),
    .B2(_14890_),
    .ZN(_11794_));
 OAI21_X1 _21138_ (.A(_11794_),
    .B1(_11401_),
    .B2(_11312_),
    .ZN(_11795_));
 OAI221_X2 _21139_ (.A(_11291_),
    .B1(_11236_),
    .B2(_11442_),
    .C1(_11428_),
    .C2(_14899_),
    .ZN(_11796_));
 NAND2_X1 _21140_ (.A1(_14899_),
    .A2(_11378_),
    .ZN(_11797_));
 AOI21_X1 _21141_ (.A(net196),
    .B1(_11382_),
    .B2(_11797_),
    .ZN(_11798_));
 OAI22_X2 _21142_ (.A1(_11292_),
    .A2(_11795_),
    .B1(_11796_),
    .B2(_11798_),
    .ZN(_11799_));
 OAI33_X1 _21143_ (.A1(_11789_),
    .A2(_11792_),
    .A3(_11793_),
    .B1(_11799_),
    .B2(_11298_),
    .B3(_11212_),
    .ZN(_11800_));
 NAND2_X1 _21144_ (.A1(_14896_),
    .A2(_11414_),
    .ZN(_11801_));
 MUX2_X1 _21145_ (.A(_11214_),
    .B(_11134_),
    .S(_11332_),
    .Z(_11802_));
 OAI221_X1 _21146_ (.A(_11405_),
    .B1(_11279_),
    .B2(_11801_),
    .C1(_11802_),
    .C2(_11330_),
    .ZN(_11803_));
 NAND4_X1 _21147_ (.A1(_11283_),
    .A2(_11178_),
    .A3(_11346_),
    .A4(_11347_),
    .ZN(_11804_));
 OAI21_X1 _21148_ (.A(_11804_),
    .B1(_11414_),
    .B2(_14904_),
    .ZN(_11805_));
 NAND2_X1 _21149_ (.A1(_11298_),
    .A2(_11805_),
    .ZN(_11806_));
 NAND3_X1 _21150_ (.A1(_11292_),
    .A2(_11803_),
    .A3(_11806_),
    .ZN(_11807_));
 MUX2_X1 _21151_ (.A(_11402_),
    .B(_11368_),
    .S(_11181_),
    .Z(_11808_));
 MUX2_X1 _21152_ (.A(_14918_),
    .B(_11808_),
    .S(_11304_),
    .Z(_11809_));
 NAND2_X2 _21153_ (.A1(_11809_),
    .A2(_11298_),
    .ZN(_11810_));
 NAND2_X1 _21154_ (.A1(_11405_),
    .A2(_11458_),
    .ZN(_11811_));
 OAI221_X2 _21155_ (.A(_14908_),
    .B1(_11295_),
    .B2(_11257_),
    .C1(_11543_),
    .C2(_11577_),
    .ZN(_11812_));
 NAND4_X4 _21156_ (.A1(_11810_),
    .A2(_11300_),
    .A3(_11811_),
    .A4(_11812_),
    .ZN(_11813_));
 AOI21_X4 _21157_ (.A(_11563_),
    .B1(_11813_),
    .B2(_11807_),
    .ZN(_11814_));
 AOI21_X1 _21158_ (.A(_11178_),
    .B1(_11323_),
    .B2(_11447_),
    .ZN(_11815_));
 AOI21_X1 _21159_ (.A(_11815_),
    .B1(_11526_),
    .B2(_11333_),
    .ZN(_11816_));
 NOR3_X2 _21160_ (.A1(_11194_),
    .A2(_11292_),
    .A3(_11816_),
    .ZN(_11817_));
 AND2_X1 _21161_ (.A1(_11331_),
    .A2(_11394_),
    .ZN(_11818_));
 AOI221_X2 _21162_ (.A(_11317_),
    .B1(_11396_),
    .B2(_11818_),
    .C1(_11484_),
    .C2(_11182_),
    .ZN(_11819_));
 NOR2_X1 _21163_ (.A1(_11322_),
    .A2(_11178_),
    .ZN(_11820_));
 AOI211_X2 _21164_ (.A(_11181_),
    .B(_11455_),
    .C1(_11373_),
    .C2(_11133_),
    .ZN(_11821_));
 NOR3_X1 _21165_ (.A1(_11291_),
    .A2(_11820_),
    .A3(_11821_),
    .ZN(_11822_));
 NOR3_X1 _21166_ (.A1(_11388_),
    .A2(_11819_),
    .A3(_11822_),
    .ZN(_11823_));
 OAI221_X2 _21167_ (.A(_11600_),
    .B1(_11678_),
    .B2(_11333_),
    .C1(_11647_),
    .C2(_11368_),
    .ZN(_11824_));
 NAND3_X1 _21168_ (.A1(_11358_),
    .A2(_11298_),
    .A3(_11824_),
    .ZN(_11825_));
 NOR3_X2 _21169_ (.A1(_11817_),
    .A2(_11823_),
    .A3(_11825_),
    .ZN(_11826_));
 OAI22_X1 _21170_ (.A1(_11155_),
    .A2(_11236_),
    .B1(_11494_),
    .B2(_11373_),
    .ZN(_11827_));
 AOI221_X2 _21171_ (.A(_11296_),
    .B1(_11400_),
    .B2(net734),
    .C1(_11827_),
    .C2(_11133_),
    .ZN(_11828_));
 AND3_X1 _21172_ (.A1(_11337_),
    .A2(_11454_),
    .A3(_11596_),
    .ZN(_11829_));
 OR3_X1 _21173_ (.A1(_11719_),
    .A2(_11828_),
    .A3(_11829_),
    .ZN(_11830_));
 AOI21_X1 _21174_ (.A(_11378_),
    .B1(_11279_),
    .B2(_11330_),
    .ZN(_11831_));
 NOR2_X1 _21175_ (.A1(net197),
    .A2(_11831_),
    .ZN(_11832_));
 NOR3_X1 _21176_ (.A1(_14896_),
    .A2(_11400_),
    .A3(_11361_),
    .ZN(_11833_));
 OAI21_X1 _21177_ (.A(_11329_),
    .B1(_11432_),
    .B2(_11833_),
    .ZN(_11834_));
 OAI21_X1 _21178_ (.A(_11439_),
    .B1(_11236_),
    .B2(_14899_),
    .ZN(_11835_));
 NAND2_X1 _21179_ (.A1(_11437_),
    .A2(_11835_),
    .ZN(_11836_));
 NAND4_X1 _21180_ (.A1(_11292_),
    .A2(_11639_),
    .A3(_11834_),
    .A4(_11836_),
    .ZN(_11837_));
 OAI21_X1 _21181_ (.A(_11830_),
    .B1(_11832_),
    .B2(_11837_),
    .ZN(_11838_));
 NOR4_X4 _21182_ (.A1(_11814_),
    .A2(_11800_),
    .A3(_11826_),
    .A4(_11838_),
    .ZN(_00063_));
 INV_X1 _21183_ (.A(_06255_),
    .ZN(_11839_));
 NOR2_X1 _21184_ (.A1(_11839_),
    .A2(_09102_),
    .ZN(_11840_));
 BUF_X8 _21185_ (.A(_08993_),
    .Z(_11841_));
 NOR2_X1 _21186_ (.A1(_06255_),
    .A2(_11841_),
    .ZN(_11842_));
 XNOR2_X2 _21187_ (.A(_08979_),
    .B(_09151_),
    .ZN(_11843_));
 XNOR2_X2 _21188_ (.A(\sa00_sr[1] ),
    .B(_08987_),
    .ZN(_11844_));
 XNOR2_X2 _21189_ (.A(_11843_),
    .B(_11844_),
    .ZN(_11845_));
 XNOR2_X1 _21190_ (.A(\sa20_sr[1] ),
    .B(_09007_),
    .ZN(_11846_));
 XNOR2_X2 _21191_ (.A(_11845_),
    .B(_11846_),
    .ZN(_11847_));
 MUX2_X2 _21192_ (.A(_11840_),
    .B(_11842_),
    .S(_11847_),
    .Z(_11848_));
 NAND3_X2 _21193_ (.A1(_06255_),
    .A2(_09728_),
    .A3(_00452_),
    .ZN(_11849_));
 NAND2_X1 _21194_ (.A1(_11839_),
    .A2(_08974_),
    .ZN(_11850_));
 OAI21_X4 _21195_ (.A(_11849_),
    .B1(_11850_),
    .B2(_00452_),
    .ZN(_11851_));
 NOR2_X4 _21196_ (.A1(_11851_),
    .A2(_11848_),
    .ZN(_11852_));
 INV_X8 _21197_ (.A(net841),
    .ZN(_11853_));
 BUF_X4 clone109 (.A(_11852_),
    .Z(net109));
 BUF_X16 _21199_ (.A(_11853_),
    .Z(_11855_));
 BUF_X32 _21200_ (.A(_11855_),
    .Z(_14928_));
 XNOR2_X2 _21201_ (.A(\sa00_sr[0] ),
    .B(\sa30_sr[0] ),
    .ZN(_11856_));
 XNOR2_X1 _21202_ (.A(net1102),
    .B(net692),
    .ZN(_11857_));
 XOR2_X2 _21203_ (.A(_08979_),
    .B(_09151_),
    .Z(_11858_));
 NAND3_X1 _21204_ (.A1(_06241_),
    .A2(_09011_),
    .A3(_11858_),
    .ZN(_11859_));
 NOR2_X1 _21205_ (.A1(_06241_),
    .A2(_08992_),
    .ZN(_11860_));
 NAND2_X1 _21206_ (.A1(net840),
    .A2(_11860_),
    .ZN(_11861_));
 AOI21_X1 _21207_ (.A(_11857_),
    .B1(_11859_),
    .B2(_11861_),
    .ZN(_11862_));
 XOR2_X1 _21208_ (.A(net692),
    .B(net1102),
    .Z(_11863_));
 NAND2_X1 _21209_ (.A1(_11858_),
    .A2(_11860_),
    .ZN(_11864_));
 NAND3_X1 _21210_ (.A1(_06241_),
    .A2(_09022_),
    .A3(net840),
    .ZN(_11865_));
 AOI21_X1 _21211_ (.A(_11863_),
    .B1(_11864_),
    .B2(_11865_),
    .ZN(_11866_));
 INV_X1 _21212_ (.A(_06241_),
    .ZN(_11867_));
 NAND3_X1 _21213_ (.A1(_11867_),
    .A2(_09726_),
    .A3(_00453_),
    .ZN(_11868_));
 NAND2_X1 _21214_ (.A1(_06241_),
    .A2(_09027_),
    .ZN(_11869_));
 OAI21_X1 _21215_ (.A(_11868_),
    .B1(_11869_),
    .B2(_00453_),
    .ZN(_11870_));
 OR3_X4 _21216_ (.A1(_11866_),
    .A2(_11862_),
    .A3(_11870_),
    .ZN(_11871_));
 BUF_X16 _21217_ (.A(_11871_),
    .Z(_11872_));
 INV_X4 _21218_ (.A(_11872_),
    .ZN(_11873_));
 BUF_X16 _21219_ (.A(_11873_),
    .Z(_11874_));
 BUF_X8 _21220_ (.A(_11874_),
    .Z(_14931_));
 XNOR2_X2 _21221_ (.A(_09037_),
    .B(_09088_),
    .ZN(_11875_));
 XNOR2_X1 _21222_ (.A(_09041_),
    .B(_11875_),
    .ZN(_11876_));
 XOR2_X2 _21223_ (.A(net629),
    .B(net695),
    .Z(_11877_));
 NAND3_X1 _21224_ (.A1(_06296_),
    .A2(_09074_),
    .A3(_11877_),
    .ZN(_11878_));
 NOR2_X1 _21225_ (.A1(net1003),
    .A2(_08972_),
    .ZN(_11879_));
 NAND2_X1 _21226_ (.A1(net922),
    .A2(_11879_),
    .ZN(_11880_));
 AOI21_X2 _21227_ (.A(_11876_),
    .B1(_11878_),
    .B2(_11880_),
    .ZN(_11881_));
 XOR2_X2 _21228_ (.A(_09037_),
    .B(_09088_),
    .Z(_11882_));
 XNOR2_X1 _21229_ (.A(_09041_),
    .B(_11882_),
    .ZN(_11883_));
 NAND2_X1 _21230_ (.A1(_11877_),
    .A2(_11879_),
    .ZN(_11884_));
 NAND3_X1 _21231_ (.A1(_06296_),
    .A2(_09011_),
    .A3(net922),
    .ZN(_11885_));
 AOI21_X2 _21232_ (.A(_11883_),
    .B1(_11884_),
    .B2(_11885_),
    .ZN(_11886_));
 INV_X1 _21233_ (.A(net1003),
    .ZN(_11887_));
 NAND3_X1 _21234_ (.A1(_11887_),
    .A2(_08993_),
    .A3(_00454_),
    .ZN(_11888_));
 NAND2_X1 _21235_ (.A1(_06296_),
    .A2(_08993_),
    .ZN(_11889_));
 OAI21_X2 _21236_ (.A(_11888_),
    .B1(_11889_),
    .B2(_00454_),
    .ZN(_11890_));
 NOR3_X4 _21237_ (.A1(_11881_),
    .A2(_11886_),
    .A3(_11890_),
    .ZN(_11891_));
 INV_X4 _21238_ (.A(_11891_),
    .ZN(_11892_));
 BUF_X4 _21239_ (.A(_11892_),
    .Z(_11893_));
 BUF_X4 _21240_ (.A(_11893_),
    .Z(_11894_));
 BUF_X4 _21241_ (.A(_11894_),
    .Z(_14947_));
 BUF_X8 _21242_ (.A(_11872_),
    .Z(_14922_));
 BUF_X4 _21243_ (.A(_11891_),
    .Z(_11895_));
 BUF_X4 _21244_ (.A(_11895_),
    .Z(_11896_));
 BUF_X4 _21245_ (.A(_11896_),
    .Z(_14940_));
 XNOR2_X2 _21246_ (.A(_09071_),
    .B(_09154_),
    .ZN(_11897_));
 XNOR2_X1 _21247_ (.A(_09165_),
    .B(_09067_),
    .ZN(_11898_));
 XNOR2_X1 _21248_ (.A(_11897_),
    .B(_11898_),
    .ZN(_11899_));
 XNOR2_X1 _21249_ (.A(_09070_),
    .B(_11899_),
    .ZN(_11900_));
 MUX2_X2 _21250_ (.A(\text_in_r[118] ),
    .B(_11900_),
    .S(_10571_),
    .Z(_11901_));
 XNOR2_X2 _21251_ (.A(_06575_),
    .B(_11901_),
    .ZN(_11902_));
 BUF_X4 _21252_ (.A(_11902_),
    .Z(_11903_));
 BUF_X4 _21253_ (.A(_11903_),
    .Z(_11904_));
 BUF_X4 _21254_ (.A(_11904_),
    .Z(_11905_));
 XNOR2_X1 _21255_ (.A(_09190_),
    .B(_09151_),
    .ZN(_11906_));
 XNOR2_X2 _21256_ (.A(_09089_),
    .B(_11906_),
    .ZN(_11907_));
 XOR2_X1 _21257_ (.A(_09187_),
    .B(_09162_),
    .Z(_11908_));
 XNOR2_X1 _21258_ (.A(_09093_),
    .B(_11908_),
    .ZN(_11909_));
 XNOR2_X1 _21259_ (.A(_11907_),
    .B(_11909_),
    .ZN(_11910_));
 MUX2_X2 _21260_ (.A(\text_in_r[116] ),
    .B(_11910_),
    .S(_09116_),
    .Z(_11911_));
 XOR2_X2 _21261_ (.A(_06281_),
    .B(_11911_),
    .Z(_11912_));
 BUF_X4 _21262_ (.A(_11912_),
    .Z(_11913_));
 CLKBUF_X3 _21263_ (.A(_11913_),
    .Z(_11914_));
 CLKBUF_X3 _21264_ (.A(_14924_),
    .Z(_11915_));
 INV_X4 _21265_ (.A(_11915_),
    .ZN(_11916_));
 NAND2_X1 _21266_ (.A1(_06221_),
    .A2(net949),
    .ZN(_11917_));
 INV_X1 _21267_ (.A(_06221_),
    .ZN(_11918_));
 NAND2_X1 _21268_ (.A1(_11918_),
    .A2(net949),
    .ZN(_11919_));
 XNOR2_X1 _21269_ (.A(_09042_),
    .B(net1101),
    .ZN(_11920_));
 XOR2_X2 _21270_ (.A(_09094_),
    .B(_09186_),
    .Z(_11921_));
 XNOR2_X2 _21271_ (.A(_09089_),
    .B(_11921_),
    .ZN(_11922_));
 XNOR2_X2 _21272_ (.A(_11920_),
    .B(_11922_),
    .ZN(_11923_));
 MUX2_X1 _21273_ (.A(_11917_),
    .B(_11919_),
    .S(_11923_),
    .Z(_11924_));
 BUF_X8 _21274_ (.A(_11924_),
    .Z(_11925_));
 BUF_X4 _21275_ (.A(_11925_),
    .Z(_11926_));
 OR3_X2 _21276_ (.A1(_11918_),
    .A2(_09099_),
    .A3(\text_in_r[115] ),
    .ZN(_11927_));
 NAND3_X2 _21277_ (.A1(_11918_),
    .A2(_09102_),
    .A3(\text_in_r[115] ),
    .ZN(_11928_));
 AND2_X1 _21278_ (.A1(_11927_),
    .A2(_11928_),
    .ZN(_11929_));
 BUF_X8 _21279_ (.A(_11929_),
    .Z(_11930_));
 BUF_X4 _21280_ (.A(_11930_),
    .Z(_11931_));
 NAND3_X2 _21281_ (.A1(_11892_),
    .A2(_11926_),
    .A3(_11931_),
    .ZN(_11932_));
 BUF_X4 _21282_ (.A(_11932_),
    .Z(_11933_));
 NOR2_X1 _21283_ (.A1(_11916_),
    .A2(_11933_),
    .ZN(_11934_));
 BUF_X2 clone110 (.A(net111),
    .Z(net110));
 NAND3_X2 _21285_ (.A1(_11931_),
    .A2(_11926_),
    .A3(_14926_),
    .ZN(_11936_));
 BUF_X16 _21286_ (.A(net979),
    .Z(_11937_));
 BUF_X8 _21287_ (.A(_08993_),
    .Z(_11938_));
 NOR2_X1 _21288_ (.A1(_11918_),
    .A2(_11938_),
    .ZN(_11939_));
 NOR2_X1 _21289_ (.A1(_06221_),
    .A2(_11938_),
    .ZN(_11940_));
 MUX2_X1 _21290_ (.A(_11939_),
    .B(_11940_),
    .S(_11923_),
    .Z(_11941_));
 BUF_X8 _21291_ (.A(_11941_),
    .Z(_11942_));
 BUF_X4 _21292_ (.A(_11942_),
    .Z(_11943_));
 NAND2_X4 _21293_ (.A1(_11927_),
    .A2(_11928_),
    .ZN(_11944_));
 BUF_X4 _21294_ (.A(_11944_),
    .Z(_11945_));
 OAI21_X4 _21295_ (.A(_11937_),
    .B1(_11943_),
    .B2(_11945_),
    .ZN(_11946_));
 AND3_X4 _21296_ (.A1(_11896_),
    .A2(_11936_),
    .A3(_11946_),
    .ZN(_11947_));
 OAI21_X2 _21297_ (.A(_11914_),
    .B1(_11934_),
    .B2(_11947_),
    .ZN(_11948_));
 XNOR2_X1 _21298_ (.A(_09161_),
    .B(_09065_),
    .ZN(_11949_));
 XNOR2_X2 _21299_ (.A(_09187_),
    .B(_11949_),
    .ZN(_11950_));
 NAND3_X2 _21300_ (.A1(_06269_),
    .A2(_11192_),
    .A3(_09167_),
    .ZN(_11951_));
 NOR2_X1 _21301_ (.A1(_06269_),
    .A2(_09823_),
    .ZN(_11952_));
 NAND2_X1 _21302_ (.A1(_09169_),
    .A2(_11952_),
    .ZN(_11953_));
 AOI21_X4 _21303_ (.A(_11950_),
    .B1(_11951_),
    .B2(_11953_),
    .ZN(_11954_));
 NAND3_X1 _21304_ (.A1(_09167_),
    .A2(_11950_),
    .A3(_11952_),
    .ZN(_11955_));
 NAND4_X1 _21305_ (.A1(_06269_),
    .A2(_11192_),
    .A3(_09169_),
    .A4(_11950_),
    .ZN(_11956_));
 NAND2_X2 _21306_ (.A1(_11955_),
    .A2(_11956_),
    .ZN(_11957_));
 OR3_X1 _21307_ (.A1(_06269_),
    .A2(_11191_),
    .A3(\text_in_r[117] ),
    .ZN(_11958_));
 NAND3_X1 _21308_ (.A1(_06269_),
    .A2(_08996_),
    .A3(\text_in_r[117] ),
    .ZN(_11959_));
 NAND2_X2 _21309_ (.A1(_11958_),
    .A2(_11959_),
    .ZN(_11960_));
 OR3_X4 _21310_ (.A1(_11954_),
    .A2(_11957_),
    .A3(_11960_),
    .ZN(_11961_));
 BUF_X4 _21311_ (.A(_11961_),
    .Z(_11962_));
 BUF_X4 _21312_ (.A(_11962_),
    .Z(_11963_));
 BUF_X4 _21313_ (.A(_11912_),
    .Z(_11964_));
 BUF_X4 _21314_ (.A(_11895_),
    .Z(_11965_));
 NAND2_X1 _21315_ (.A1(_11855_),
    .A2(_11965_),
    .ZN(_11966_));
 NAND2_X4 _21316_ (.A1(_11925_),
    .A2(_11930_),
    .ZN(_11967_));
 CLKBUF_X3 _21317_ (.A(_11967_),
    .Z(_11968_));
 BUF_X4 _21318_ (.A(_14925_),
    .Z(_11969_));
 INV_X8 _21319_ (.A(_11969_),
    .ZN(_11970_));
 NOR2_X4 _21320_ (.A1(_11970_),
    .A2(_11891_),
    .ZN(_11971_));
 NOR2_X2 _21321_ (.A1(_11968_),
    .A2(_11971_),
    .ZN(_11972_));
 AOI21_X4 _21322_ (.A(_11964_),
    .B1(_11972_),
    .B2(_11966_),
    .ZN(_11973_));
 BUF_X4 _21323_ (.A(_11967_),
    .Z(_11974_));
 BUF_X4 _21324_ (.A(_11974_),
    .Z(_11975_));
 BUF_X4 _21325_ (.A(_14932_),
    .Z(_11976_));
 NOR2_X1 _21326_ (.A1(_11976_),
    .A2(_11965_),
    .ZN(_11977_));
 NOR2_X2 _21327_ (.A1(_11872_),
    .A2(_11892_),
    .ZN(_11978_));
 CLKBUF_X3 _21328_ (.A(_11978_),
    .Z(_11979_));
 OAI21_X1 _21329_ (.A(_11975_),
    .B1(_11977_),
    .B2(_11979_),
    .ZN(_11980_));
 AOI21_X2 _21330_ (.A(_11963_),
    .B1(_11980_),
    .B2(_11973_),
    .ZN(_11981_));
 AOI21_X4 _21331_ (.A(_11891_),
    .B1(_11926_),
    .B2(_11931_),
    .ZN(_11982_));
 NOR2_X4 _21332_ (.A1(_11874_),
    .A2(_11891_),
    .ZN(_11983_));
 AOI221_X2 _21333_ (.A(_11983_),
    .B1(_11931_),
    .B2(_11926_),
    .C1(_11853_),
    .C2(_11978_),
    .ZN(_11984_));
 OAI21_X1 _21334_ (.A(_11982_),
    .B1(_11984_),
    .B2(_11964_),
    .ZN(_11985_));
 XNOR2_X2 _21335_ (.A(_06281_),
    .B(_11911_),
    .ZN(_11986_));
 BUF_X4 _21336_ (.A(_11986_),
    .Z(_11987_));
 BUF_X4 _21337_ (.A(_11987_),
    .Z(_11988_));
 BUF_X4 _21338_ (.A(_11892_),
    .Z(_11989_));
 BUF_X4 _21339_ (.A(_11989_),
    .Z(_11990_));
 NAND3_X4 _21340_ (.A1(_14934_),
    .A2(_11925_),
    .A3(_11930_),
    .ZN(_11991_));
 OAI21_X1 _21341_ (.A(net1199),
    .B1(_11943_),
    .B2(_11945_),
    .ZN(_11992_));
 AOI21_X1 _21342_ (.A(_11990_),
    .B1(_11991_),
    .B2(_11992_),
    .ZN(_11993_));
 NOR2_X1 _21343_ (.A1(_11988_),
    .A2(_11993_),
    .ZN(_11994_));
 NOR2_X2 _21344_ (.A1(_11913_),
    .A2(_11984_),
    .ZN(_11995_));
 INV_X8 _21345_ (.A(_11937_),
    .ZN(_11996_));
 OAI221_X2 _21346_ (.A(_11985_),
    .B1(_11994_),
    .B2(_11995_),
    .C1(_11996_),
    .C2(_11933_),
    .ZN(_11997_));
 BUF_X4 _21347_ (.A(_11963_),
    .Z(_11998_));
 AOI221_X2 _21348_ (.A(_11905_),
    .B1(_11948_),
    .B2(_11981_),
    .C1(_11997_),
    .C2(_11998_),
    .ZN(_11999_));
 XOR2_X1 _21349_ (.A(_09068_),
    .B(net609),
    .Z(_12000_));
 XNOR2_X1 _21350_ (.A(_08978_),
    .B(_12000_),
    .ZN(_12001_));
 MUX2_X2 _21351_ (.A(\text_in_r[119] ),
    .B(_12001_),
    .S(_09076_),
    .Z(_12002_));
 XOR2_X2 _21352_ (.A(_06587_),
    .B(_12002_),
    .Z(_12003_));
 CLKBUF_X3 _21353_ (.A(_12003_),
    .Z(_12004_));
 NOR3_X4 _21354_ (.A1(_11954_),
    .A2(_11957_),
    .A3(_11960_),
    .ZN(_12005_));
 CLKBUF_X3 _21355_ (.A(_12005_),
    .Z(_12006_));
 CLKBUF_X3 _21356_ (.A(_12006_),
    .Z(_12007_));
 CLKBUF_X3 _21357_ (.A(_11987_),
    .Z(_12008_));
 CLKBUF_X3 _21358_ (.A(_11968_),
    .Z(_12009_));
 NOR3_X4 _21359_ (.A1(_11891_),
    .A2(_11942_),
    .A3(_11944_),
    .ZN(_12010_));
 CLKBUF_X3 _21360_ (.A(_11969_),
    .Z(_12011_));
 AOI22_X1 _21361_ (.A1(_14945_),
    .A2(_12009_),
    .B1(_12010_),
    .B2(_12011_),
    .ZN(_12012_));
 OR2_X1 _21362_ (.A1(_12008_),
    .A2(_12012_),
    .ZN(_12013_));
 CLKBUF_X3 _21363_ (.A(_11988_),
    .Z(_12014_));
 NOR2_X4 _21364_ (.A1(_11874_),
    .A2(_11892_),
    .ZN(_12015_));
 BUF_X4 _21365_ (.A(_11853_),
    .Z(_12016_));
 NOR2_X4 _21366_ (.A1(_14929_),
    .A2(_14926_),
    .ZN(_12017_));
 AOI221_X2 _21367_ (.A(_11968_),
    .B1(_12015_),
    .B2(_12016_),
    .C1(net1098),
    .C2(_11894_),
    .ZN(_12018_));
 NOR2_X4 _21368_ (.A1(_11942_),
    .A2(_11944_),
    .ZN(_12019_));
 BUF_X4 _21369_ (.A(_12019_),
    .Z(_12020_));
 CLKBUF_X3 _21370_ (.A(_12020_),
    .Z(_12021_));
 CLKBUF_X3 _21371_ (.A(_12021_),
    .Z(_12022_));
 BUF_X4 _21372_ (.A(_11965_),
    .Z(_12023_));
 NAND2_X1 _21373_ (.A1(_11916_),
    .A2(_12023_),
    .ZN(_12024_));
 NAND2_X1 _21374_ (.A1(_14931_),
    .A2(_11894_),
    .ZN(_12025_));
 AOI21_X1 _21375_ (.A(_12022_),
    .B1(_12024_),
    .B2(_12025_),
    .ZN(_12026_));
 OAI21_X1 _21376_ (.A(_12014_),
    .B1(_12018_),
    .B2(_12026_),
    .ZN(_12027_));
 AOI21_X1 _21377_ (.A(_12007_),
    .B1(_12013_),
    .B2(_12027_),
    .ZN(_12028_));
 BUF_X8 _21378_ (.A(_14934_),
    .Z(_12029_));
 INV_X4 _21379_ (.A(net1200),
    .ZN(_12030_));
 BUF_X4 _21380_ (.A(_12019_),
    .Z(_12031_));
 AOI21_X4 _21381_ (.A(_11874_),
    .B1(_11925_),
    .B2(_11930_),
    .ZN(_12032_));
 AOI22_X2 _21382_ (.A1(_12030_),
    .A2(_12031_),
    .B1(_12032_),
    .B2(_12016_),
    .ZN(_12033_));
 AOI221_X2 _21383_ (.A(_11964_),
    .B1(_11982_),
    .B2(_12029_),
    .C1(_12033_),
    .C2(_12023_),
    .ZN(_12034_));
 OAI21_X2 _21384_ (.A(_11895_),
    .B1(_11943_),
    .B2(_11945_),
    .ZN(_12035_));
 OAI21_X4 _21385_ (.A(_11912_),
    .B1(_12030_),
    .B2(_12035_),
    .ZN(_12036_));
 AOI221_X1 _21386_ (.A(_11968_),
    .B1(_12015_),
    .B2(_12016_),
    .C1(_11894_),
    .C2(_11976_),
    .ZN(_12037_));
 OAI21_X1 _21387_ (.A(_12006_),
    .B1(_12036_),
    .B2(_12037_),
    .ZN(_12038_));
 OAI21_X1 _21388_ (.A(_11905_),
    .B1(_12034_),
    .B2(_12038_),
    .ZN(_12039_));
 OAI21_X1 _21389_ (.A(_12004_),
    .B1(_12028_),
    .B2(_12039_),
    .ZN(_12040_));
 BUF_X4 _21390_ (.A(_11964_),
    .Z(_12041_));
 NAND3_X2 _21391_ (.A1(_11969_),
    .A2(_11926_),
    .A3(_11931_),
    .ZN(_12042_));
 CLKBUF_X3 _21392_ (.A(_11895_),
    .Z(_12043_));
 NOR2_X1 _21393_ (.A1(_12016_),
    .A2(_12043_),
    .ZN(_12044_));
 NAND2_X4 _21394_ (.A1(_11970_),
    .A2(_11989_),
    .ZN(_12045_));
 NOR2_X2 _21395_ (.A1(_12016_),
    .A2(_11968_),
    .ZN(_12046_));
 OAI221_X2 _21396_ (.A(_11904_),
    .B1(_12042_),
    .B2(_12044_),
    .C1(_12045_),
    .C2(_12046_),
    .ZN(_12047_));
 BUF_X2 rebuffer635 (.A(net1099),
    .Z(net1098));
 INV_X2 _21398_ (.A(_14938_),
    .ZN(_12049_));
 AOI21_X4 _21399_ (.A(_12049_),
    .B1(_11926_),
    .B2(_11931_),
    .ZN(_12050_));
 AOI21_X1 _21400_ (.A(_12050_),
    .B1(_12021_),
    .B2(_14928_),
    .ZN(_12051_));
 BUF_X8 _21401_ (.A(_11852_),
    .Z(_12052_));
 NAND2_X2 _21402_ (.A1(_12052_),
    .A2(_12031_),
    .ZN(_12053_));
 AOI22_X1 _21403_ (.A1(_14940_),
    .A2(_12051_),
    .B1(_12053_),
    .B2(_11983_),
    .ZN(_12054_));
 OAI21_X1 _21404_ (.A(_12047_),
    .B1(_12054_),
    .B2(_11905_),
    .ZN(_12055_));
 AND2_X1 _21405_ (.A1(_12041_),
    .A2(_12055_),
    .ZN(_12056_));
 NOR2_X1 _21406_ (.A1(_12006_),
    .A2(_12003_),
    .ZN(_12057_));
 XOR2_X2 _21407_ (.A(_06575_),
    .B(_11901_),
    .Z(_12058_));
 BUF_X4 _21408_ (.A(_12058_),
    .Z(_12059_));
 NOR2_X2 _21409_ (.A1(_11914_),
    .A2(_12059_),
    .ZN(_12060_));
 NOR3_X4 _21410_ (.A1(_11892_),
    .A2(_11942_),
    .A3(_11944_),
    .ZN(_12061_));
 NOR2_X4 _21411_ (.A1(_11982_),
    .A2(_12061_),
    .ZN(_12062_));
 NOR2_X1 _21412_ (.A1(_11916_),
    .A2(_12062_),
    .ZN(_12063_));
 INV_X2 _21413_ (.A(_11976_),
    .ZN(_12064_));
 CLKBUF_X3 _21414_ (.A(_12035_),
    .Z(_12065_));
 OAI22_X1 _21415_ (.A1(_12064_),
    .A2(_11933_),
    .B1(_12065_),
    .B2(_12011_),
    .ZN(_12066_));
 OAI21_X1 _21416_ (.A(_12060_),
    .B1(_12063_),
    .B2(_12066_),
    .ZN(_12067_));
 BUF_X16 _21417_ (.A(_12052_),
    .Z(_12068_));
 BUF_X4 _21418_ (.A(_11990_),
    .Z(_12069_));
 MUX2_X1 _21419_ (.A(_14926_),
    .B(net715),
    .S(_12069_),
    .Z(_12070_));
 AOI21_X1 _21420_ (.A(_11905_),
    .B1(_12070_),
    .B2(_12022_),
    .ZN(_12071_));
 NAND2_X1 _21421_ (.A1(_11995_),
    .A2(_12071_),
    .ZN(_12072_));
 NAND3_X1 _21422_ (.A1(_12057_),
    .A2(_12067_),
    .A3(_12072_),
    .ZN(_12073_));
 XNOR2_X2 _21423_ (.A(_06587_),
    .B(_12002_),
    .ZN(_12074_));
 BUF_X4 _21424_ (.A(_12074_),
    .Z(_12075_));
 NOR2_X2 _21425_ (.A1(_11987_),
    .A2(_12058_),
    .ZN(_12076_));
 AOI21_X1 _21426_ (.A(_11979_),
    .B1(_14922_),
    .B2(_12068_),
    .ZN(_12077_));
 XNOR2_X1 _21427_ (.A(_12009_),
    .B(_12077_),
    .ZN(_12078_));
 NAND2_X1 _21428_ (.A1(_12076_),
    .A2(_12078_),
    .ZN(_12079_));
 BUF_X4 _21429_ (.A(_11990_),
    .Z(_12080_));
 OAI21_X1 _21430_ (.A(_12080_),
    .B1(_12050_),
    .B2(_12046_),
    .ZN(_12081_));
 AOI21_X4 _21431_ (.A(_11892_),
    .B1(_11925_),
    .B2(_11930_),
    .ZN(_12082_));
 NAND2_X1 _21432_ (.A1(_12011_),
    .A2(_12082_),
    .ZN(_12083_));
 NAND3_X4 _21433_ (.A1(_11874_),
    .A2(_11926_),
    .A3(_11931_),
    .ZN(_12084_));
 NOR2_X1 _21434_ (.A1(_11987_),
    .A2(_11903_),
    .ZN(_12085_));
 NAND4_X1 _21435_ (.A1(_12081_),
    .A2(_12083_),
    .A3(_12084_),
    .A4(_12085_),
    .ZN(_12086_));
 NAND4_X1 _21436_ (.A1(_12007_),
    .A2(_12075_),
    .A3(_12079_),
    .A4(_12086_),
    .ZN(_12087_));
 AOI21_X1 _21437_ (.A(_11893_),
    .B1(_11968_),
    .B2(_11976_),
    .ZN(_12088_));
 OAI21_X1 _21438_ (.A(_12088_),
    .B1(_12009_),
    .B2(_12011_),
    .ZN(_12089_));
 BUF_X8 clone213 (.A(_12052_),
    .Z(net715));
 OAI221_X1 _21440_ (.A(_14947_),
    .B1(_12021_),
    .B2(_11916_),
    .C1(_12084_),
    .C2(net715),
    .ZN(_12090_));
 AOI21_X1 _21441_ (.A(_12059_),
    .B1(_12089_),
    .B2(_12090_),
    .ZN(_12091_));
 NAND2_X2 _21442_ (.A1(net2),
    .A2(_11974_),
    .ZN(_12092_));
 AOI221_X2 _21443_ (.A(_11903_),
    .B1(_12082_),
    .B2(_11996_),
    .C1(_12092_),
    .C2(_11983_),
    .ZN(_12093_));
 NOR3_X1 _21444_ (.A1(_12041_),
    .A2(_12091_),
    .A3(_12093_),
    .ZN(_12094_));
 OAI222_X2 _21445_ (.A1(_11999_),
    .A2(_12040_),
    .B1(_12056_),
    .B2(_12073_),
    .C1(_12087_),
    .C2(_12094_),
    .ZN(_00064_));
 NAND2_X1 _21446_ (.A1(_11913_),
    .A2(_11902_),
    .ZN(_12095_));
 NOR3_X1 _21447_ (.A1(_12069_),
    .A2(_12005_),
    .A3(_12095_),
    .ZN(_12096_));
 OAI21_X1 _21448_ (.A(_12084_),
    .B1(_12020_),
    .B2(_11937_),
    .ZN(_12097_));
 AOI221_X2 _21449_ (.A(_11967_),
    .B1(_11978_),
    .B2(_11853_),
    .C1(_14932_),
    .C2(_11893_),
    .ZN(_12098_));
 INV_X1 _21450_ (.A(_12098_),
    .ZN(_12099_));
 NAND2_X1 _21451_ (.A1(_11987_),
    .A2(_11903_),
    .ZN(_12100_));
 NOR2_X1 _21452_ (.A1(_12005_),
    .A2(_12031_),
    .ZN(_12101_));
 INV_X1 _21453_ (.A(_14948_),
    .ZN(_12102_));
 AOI21_X1 _21454_ (.A(_12100_),
    .B1(_12101_),
    .B2(_12102_),
    .ZN(_12103_));
 AOI221_X1 _21455_ (.A(_12003_),
    .B1(_12096_),
    .B2(_12097_),
    .C1(_12099_),
    .C2(_12103_),
    .ZN(_12104_));
 NOR2_X1 _21456_ (.A1(_11916_),
    .A2(_11895_),
    .ZN(_12105_));
 OAI21_X1 _21457_ (.A(_12022_),
    .B1(_12015_),
    .B2(_12105_),
    .ZN(_12106_));
 OAI221_X1 _21458_ (.A(_14928_),
    .B1(_11943_),
    .B2(_11945_),
    .C1(_11983_),
    .C2(_11979_),
    .ZN(_12107_));
 AOI21_X1 _21459_ (.A(_11998_),
    .B1(_12106_),
    .B2(_12107_),
    .ZN(_12108_));
 BUF_X4 _21460_ (.A(_12020_),
    .Z(_12109_));
 NAND2_X1 _21461_ (.A1(_11855_),
    .A2(_12109_),
    .ZN(_12110_));
 AOI21_X1 _21462_ (.A(_12023_),
    .B1(_12110_),
    .B2(_12092_),
    .ZN(_12111_));
 AOI21_X1 _21463_ (.A(_12108_),
    .B1(_12111_),
    .B2(_11998_),
    .ZN(_12112_));
 OAI21_X1 _21464_ (.A(_12104_),
    .B1(_12112_),
    .B2(_12095_),
    .ZN(_12113_));
 AOI21_X4 _21465_ (.A(_11969_),
    .B1(_11925_),
    .B2(_11930_),
    .ZN(_12114_));
 NOR3_X4 _21466_ (.A1(_11872_),
    .A2(_11943_),
    .A3(_11945_),
    .ZN(_12115_));
 AOI21_X1 _21467_ (.A(net1012),
    .B1(_12115_),
    .B2(_14928_),
    .ZN(_12116_));
 OAI221_X1 _21468_ (.A(_12008_),
    .B1(_11933_),
    .B2(_14931_),
    .C1(_12116_),
    .C2(_14947_),
    .ZN(_12117_));
 NAND3_X4 _21469_ (.A1(_14938_),
    .A2(_11925_),
    .A3(_11930_),
    .ZN(_12118_));
 NAND2_X1 _21470_ (.A1(_12023_),
    .A2(_12118_),
    .ZN(_12119_));
 OAI21_X4 _21471_ (.A(_11873_),
    .B1(_11851_),
    .B2(net553),
    .ZN(_12120_));
 MUX2_X1 _21472_ (.A(_14926_),
    .B(_12120_),
    .S(_11974_),
    .Z(_12121_));
 OAI221_X1 _21473_ (.A(_12041_),
    .B1(net1012),
    .B2(_12119_),
    .C1(_12121_),
    .C2(_14940_),
    .ZN(_12122_));
 AND4_X1 _21474_ (.A1(_11998_),
    .A2(_12059_),
    .A3(_12117_),
    .A4(_12122_),
    .ZN(_12123_));
 MUX2_X1 _21475_ (.A(_11915_),
    .B(net2),
    .S(_11967_),
    .Z(_12124_));
 MUX2_X1 _21476_ (.A(_12097_),
    .B(_12124_),
    .S(_11894_),
    .Z(_12125_));
 OR2_X1 _21477_ (.A1(_12041_),
    .A2(_12125_),
    .ZN(_12126_));
 AOI21_X4 _21478_ (.A(_11970_),
    .B1(_11926_),
    .B2(_11931_),
    .ZN(_12127_));
 NOR3_X4 _21479_ (.A1(_12127_),
    .A2(_12043_),
    .A3(_12115_),
    .ZN(_12128_));
 OAI21_X2 _21480_ (.A(_11936_),
    .B1(_12031_),
    .B2(_11915_),
    .ZN(_12129_));
 NOR2_X1 _21481_ (.A1(_12069_),
    .A2(_12129_),
    .ZN(_12130_));
 OR3_X4 _21482_ (.A1(_11988_),
    .A2(_12128_),
    .A3(_12130_),
    .ZN(_12131_));
 AND4_X4 _21483_ (.A1(_12007_),
    .A2(_12059_),
    .A3(_12126_),
    .A4(_12131_),
    .ZN(_12132_));
 OAI21_X4 _21484_ (.A(_11872_),
    .B1(_11942_),
    .B2(_11944_),
    .ZN(_12133_));
 AOI21_X1 _21485_ (.A(net109),
    .B1(_12069_),
    .B2(_12133_),
    .ZN(_12134_));
 NOR2_X2 _21486_ (.A1(_11961_),
    .A2(_11912_),
    .ZN(_12135_));
 NOR3_X4 _21487_ (.A1(_11874_),
    .A2(_11942_),
    .A3(_11944_),
    .ZN(_12136_));
 NAND2_X1 _21488_ (.A1(_12052_),
    .A2(_12136_),
    .ZN(_12137_));
 NAND3_X1 _21489_ (.A1(_12065_),
    .A2(_12135_),
    .A3(_12137_),
    .ZN(_12138_));
 OAI21_X1 _21490_ (.A(_11903_),
    .B1(_12134_),
    .B2(_12138_),
    .ZN(_12139_));
 NOR2_X2 _21491_ (.A1(_11962_),
    .A2(_11987_),
    .ZN(_12140_));
 NAND3_X1 _21492_ (.A1(_11990_),
    .A2(_12133_),
    .A3(_12084_),
    .ZN(_12141_));
 NOR3_X4 _21493_ (.A1(net977),
    .A2(_11942_),
    .A3(_11944_),
    .ZN(_12142_));
 OR2_X2 _21494_ (.A1(net1011),
    .A2(_12142_),
    .ZN(_12143_));
 OAI21_X2 _21495_ (.A(_12141_),
    .B1(_12143_),
    .B2(_12080_),
    .ZN(_12144_));
 OAI221_X1 _21496_ (.A(_11964_),
    .B1(_11932_),
    .B2(net978),
    .C1(_12062_),
    .C2(net715),
    .ZN(_12145_));
 NOR2_X1 _21497_ (.A1(_12049_),
    .A2(_11989_),
    .ZN(_12146_));
 OR3_X1 _21498_ (.A1(_12020_),
    .A2(_11971_),
    .A3(_12146_),
    .ZN(_12147_));
 NOR2_X4 _21499_ (.A1(_11937_),
    .A2(_11895_),
    .ZN(_12148_));
 AOI21_X4 _21500_ (.A(_12148_),
    .B1(_12015_),
    .B2(_12016_),
    .ZN(_12149_));
 OAI21_X1 _21501_ (.A(_12147_),
    .B1(_12149_),
    .B2(_11975_),
    .ZN(_12150_));
 OAI21_X2 _21502_ (.A(_12145_),
    .B1(_12150_),
    .B2(_11914_),
    .ZN(_12151_));
 AOI221_X2 _21503_ (.A(_12139_),
    .B1(_12140_),
    .B2(_12144_),
    .C1(_11963_),
    .C2(_12151_),
    .ZN(_12152_));
 BUF_X4 _21504_ (.A(_14938_),
    .Z(_12153_));
 OAI21_X1 _21505_ (.A(_12153_),
    .B1(_11943_),
    .B2(_11945_),
    .ZN(_12154_));
 NAND2_X1 _21506_ (.A1(_12023_),
    .A2(_12120_),
    .ZN(_12155_));
 NAND3_X1 _21507_ (.A1(_12065_),
    .A2(_12154_),
    .A3(_12155_),
    .ZN(_12156_));
 NAND2_X1 _21508_ (.A1(_12005_),
    .A2(_11913_),
    .ZN(_12157_));
 AOI21_X2 _21509_ (.A(_12157_),
    .B1(_12082_),
    .B2(net1013),
    .ZN(_12158_));
 AND2_X1 _21510_ (.A1(_12156_),
    .A2(_12158_),
    .ZN(_12159_));
 NAND2_X2 _21511_ (.A1(_12005_),
    .A2(_11986_),
    .ZN(_12160_));
 NAND2_X1 _21512_ (.A1(_12120_),
    .A2(_11967_),
    .ZN(_12161_));
 AOI21_X1 _21513_ (.A(_12114_),
    .B1(_12109_),
    .B2(net978),
    .ZN(_12162_));
 BUF_X4 _21514_ (.A(_12043_),
    .Z(_12163_));
 MUX2_X1 _21515_ (.A(_12161_),
    .B(_12162_),
    .S(_12163_),
    .Z(_12164_));
 NAND2_X1 _21516_ (.A1(_11962_),
    .A2(_11987_),
    .ZN(_12165_));
 NAND2_X1 _21517_ (.A1(net1199),
    .A2(_12010_),
    .ZN(_12166_));
 OAI21_X4 _21518_ (.A(_11874_),
    .B1(_11942_),
    .B2(_11944_),
    .ZN(_12167_));
 OAI221_X1 _21519_ (.A(_12166_),
    .B1(_12062_),
    .B2(_14931_),
    .C1(_12167_),
    .C2(_11855_),
    .ZN(_12168_));
 OAI22_X1 _21520_ (.A1(_12160_),
    .A2(_12164_),
    .B1(_12165_),
    .B2(_12168_),
    .ZN(_12169_));
 NOR3_X1 _21521_ (.A1(_11916_),
    .A2(_11943_),
    .A3(_11945_),
    .ZN(_12170_));
 OAI21_X1 _21522_ (.A(_12043_),
    .B1(_12127_),
    .B2(_12170_),
    .ZN(_12171_));
 NAND3_X1 _21523_ (.A1(_12080_),
    .A2(_11946_),
    .A3(_12084_),
    .ZN(_12172_));
 NAND4_X1 _21524_ (.A1(_11963_),
    .A2(_11914_),
    .A3(_12171_),
    .A4(_12172_),
    .ZN(_12173_));
 NAND2_X1 _21525_ (.A1(_12059_),
    .A2(_12173_),
    .ZN(_12174_));
 NOR3_X1 _21526_ (.A1(_12159_),
    .A2(_12169_),
    .A3(_12174_),
    .ZN(_12175_));
 OAI33_X1 _21527_ (.A1(_12132_),
    .A2(_12113_),
    .A3(_12123_),
    .B1(_12152_),
    .B2(_12175_),
    .B3(_12075_),
    .ZN(_00065_));
 OAI21_X4 _21528_ (.A(_12029_),
    .B1(_11943_),
    .B2(_11945_),
    .ZN(_12176_));
 NAND3_X1 _21529_ (.A1(_11896_),
    .A2(_12084_),
    .A3(_12176_),
    .ZN(_12177_));
 OAI211_X2 _21530_ (.A(_11894_),
    .B(_12118_),
    .C1(_12109_),
    .C2(_11855_),
    .ZN(_12178_));
 AOI21_X1 _21531_ (.A(_12157_),
    .B1(_12177_),
    .B2(_12178_),
    .ZN(_12179_));
 OAI211_X2 _21532_ (.A(_11896_),
    .B(_11991_),
    .C1(_12109_),
    .C2(net109),
    .ZN(_12180_));
 NOR2_X1 _21533_ (.A1(_11913_),
    .A2(_12148_),
    .ZN(_12181_));
 AOI21_X1 _21534_ (.A(_12005_),
    .B1(_12180_),
    .B2(_12181_),
    .ZN(_12182_));
 NAND3_X1 _21535_ (.A1(_11896_),
    .A2(_11991_),
    .A3(_12167_),
    .ZN(_12183_));
 NAND3_X1 _21536_ (.A1(_11990_),
    .A2(_11946_),
    .A3(_12118_),
    .ZN(_12184_));
 NAND3_X1 _21537_ (.A1(_11964_),
    .A2(_12183_),
    .A3(_12184_),
    .ZN(_12185_));
 NAND3_X1 _21538_ (.A1(_12163_),
    .A2(_11992_),
    .A3(_12084_),
    .ZN(_12186_));
 NAND2_X1 _21539_ (.A1(_12069_),
    .A2(_11991_),
    .ZN(_12187_));
 OAI21_X1 _21540_ (.A(_12186_),
    .B1(_12187_),
    .B2(net1012),
    .ZN(_12188_));
 AOI221_X2 _21541_ (.A(_12179_),
    .B1(_12182_),
    .B2(_12185_),
    .C1(_12135_),
    .C2(_12188_),
    .ZN(_12189_));
 NOR2_X1 _21542_ (.A1(_12114_),
    .A2(_12170_),
    .ZN(_12190_));
 NAND2_X1 _21543_ (.A1(_12080_),
    .A2(_12190_),
    .ZN(_12191_));
 AOI21_X1 _21544_ (.A(_12005_),
    .B1(_12053_),
    .B2(_12088_),
    .ZN(_12192_));
 NOR3_X1 _21545_ (.A1(net2),
    .A2(_12019_),
    .A3(_12015_),
    .ZN(_12193_));
 NOR2_X1 _21546_ (.A1(net1144),
    .A2(_11989_),
    .ZN(_12194_));
 MUX2_X1 _21547_ (.A(_11989_),
    .B(_12019_),
    .S(net842),
    .Z(_12195_));
 AOI221_X2 _21548_ (.A(_12193_),
    .B1(_12194_),
    .B2(_12133_),
    .C1(_11970_),
    .C2(_12195_),
    .ZN(_12196_));
 AOI221_X2 _21549_ (.A(_12008_),
    .B1(_12191_),
    .B2(_12192_),
    .C1(_12196_),
    .C2(_12006_),
    .ZN(_12197_));
 NAND3_X1 _21550_ (.A1(net1014),
    .A2(_14922_),
    .A3(_11963_),
    .ZN(_12198_));
 OR2_X1 _21551_ (.A1(_11963_),
    .A2(_12045_),
    .ZN(_12199_));
 NOR2_X1 _21552_ (.A1(_12041_),
    .A2(_12022_),
    .ZN(_12200_));
 OAI221_X1 _21553_ (.A(_14940_),
    .B1(_11962_),
    .B2(_14922_),
    .C1(_11851_),
    .C2(net555),
    .ZN(_12201_));
 NAND4_X1 _21554_ (.A1(_12198_),
    .A2(_12199_),
    .A3(_12200_),
    .A4(_12201_),
    .ZN(_12202_));
 MUX2_X1 _21555_ (.A(_14945_),
    .B(_12102_),
    .S(_11962_),
    .Z(_12203_));
 NAND3_X1 _21556_ (.A1(_12014_),
    .A2(_12022_),
    .A3(_12203_),
    .ZN(_12204_));
 NAND3_X1 _21557_ (.A1(_12004_),
    .A2(_12202_),
    .A3(_12204_),
    .ZN(_12205_));
 OAI22_X1 _21558_ (.A1(_12004_),
    .A2(_12189_),
    .B1(_12197_),
    .B2(_12205_),
    .ZN(_12206_));
 OAI221_X1 _21559_ (.A(_12135_),
    .B1(_12141_),
    .B2(net1013),
    .C1(_12153_),
    .C2(_12065_),
    .ZN(_12207_));
 NAND2_X1 _21560_ (.A1(_12074_),
    .A2(_12207_),
    .ZN(_12208_));
 NOR3_X4 _21561_ (.A1(_11942_),
    .A2(net1199),
    .A3(_11944_),
    .ZN(_12209_));
 NOR2_X1 _21562_ (.A1(_12032_),
    .A2(_12209_),
    .ZN(_12210_));
 MUX2_X1 _21563_ (.A(_14926_),
    .B(net2),
    .S(_12019_),
    .Z(_12211_));
 MUX2_X1 _21564_ (.A(_12210_),
    .B(_12211_),
    .S(_11893_),
    .Z(_12212_));
 AND2_X2 _21565_ (.A1(_12118_),
    .A2(_12167_),
    .ZN(_12213_));
 NAND2_X2 _21566_ (.A1(_11895_),
    .A2(_12020_),
    .ZN(_12214_));
 OAI221_X1 _21567_ (.A(_12092_),
    .B1(_12213_),
    .B2(_12043_),
    .C1(_12214_),
    .C2(_11996_),
    .ZN(_12215_));
 MUX2_X1 _21568_ (.A(_12212_),
    .B(_12215_),
    .S(_11962_),
    .Z(_12216_));
 NOR2_X1 _21569_ (.A1(_12021_),
    .A2(_12149_),
    .ZN(_12217_));
 NOR2_X1 _21570_ (.A1(_12006_),
    .A2(_12217_),
    .ZN(_12218_));
 AOI221_X2 _21571_ (.A(_12208_),
    .B1(_12041_),
    .B2(_12216_),
    .C1(_11973_),
    .C2(_12218_),
    .ZN(_12219_));
 AOI21_X1 _21572_ (.A(_11962_),
    .B1(_12120_),
    .B2(_11933_),
    .ZN(_12220_));
 NOR3_X1 _21573_ (.A1(_14952_),
    .A2(_12005_),
    .A3(_11975_),
    .ZN(_12221_));
 OR3_X1 _21574_ (.A1(_12008_),
    .A2(_12220_),
    .A3(_12221_),
    .ZN(_12222_));
 AOI21_X1 _21575_ (.A(_14940_),
    .B1(_11963_),
    .B2(_14922_),
    .ZN(_12223_));
 AOI21_X1 _21576_ (.A(_12223_),
    .B1(_11998_),
    .B2(net1014),
    .ZN(_12224_));
 AOI21_X1 _21577_ (.A(_12222_),
    .B1(_12224_),
    .B2(_12009_),
    .ZN(_12225_));
 AOI221_X2 _21578_ (.A(_11913_),
    .B1(_11982_),
    .B2(net978),
    .C1(_12190_),
    .C2(_12163_),
    .ZN(_12226_));
 OAI22_X1 _21579_ (.A1(_11976_),
    .A2(_11933_),
    .B1(net1098),
    .B2(_12065_),
    .ZN(_12227_));
 OAI21_X1 _21580_ (.A(_12006_),
    .B1(_12008_),
    .B2(_12227_),
    .ZN(_12228_));
 OAI21_X1 _21581_ (.A(_11872_),
    .B1(_11851_),
    .B2(net554),
    .ZN(_12229_));
 NOR3_X1 _21582_ (.A1(_14940_),
    .A2(_12009_),
    .A3(_12229_),
    .ZN(_12230_));
 NOR2_X1 _21583_ (.A1(_12006_),
    .A2(_11964_),
    .ZN(_12231_));
 INV_X1 _21584_ (.A(_14943_),
    .ZN(_12232_));
 OAI21_X1 _21585_ (.A(_12231_),
    .B1(_12022_),
    .B2(_12232_),
    .ZN(_12233_));
 OAI221_X1 _21586_ (.A(_12004_),
    .B1(_12228_),
    .B2(_12226_),
    .C1(_12230_),
    .C2(_12233_),
    .ZN(_12234_));
 OAI21_X1 _21587_ (.A(_11905_),
    .B1(_12234_),
    .B2(_12225_),
    .ZN(_12235_));
 OAI22_X2 _21588_ (.A1(_11905_),
    .A2(_12206_),
    .B1(_12219_),
    .B2(_12235_),
    .ZN(_00066_));
 AOI22_X1 _21589_ (.A1(_11979_),
    .A2(_12021_),
    .B1(_11982_),
    .B2(_14922_),
    .ZN(_12236_));
 NOR2_X1 _21590_ (.A1(net1014),
    .A2(_12236_),
    .ZN(_12237_));
 OAI221_X1 _21591_ (.A(_12008_),
    .B1(_11933_),
    .B2(_12011_),
    .C1(_12065_),
    .C2(_12064_),
    .ZN(_12238_));
 NOR2_X2 _21592_ (.A1(net842),
    .A2(_12133_),
    .ZN(_12239_));
 OAI21_X1 _21593_ (.A(_12167_),
    .B1(_11975_),
    .B2(_11976_),
    .ZN(_12240_));
 AOI221_X2 _21594_ (.A(_12239_),
    .B1(_12061_),
    .B2(_11970_),
    .C1(_12240_),
    .C2(_12080_),
    .ZN(_12241_));
 OAI221_X1 _21595_ (.A(_12007_),
    .B1(_12237_),
    .B2(_12238_),
    .C1(_12241_),
    .C2(_12014_),
    .ZN(_12242_));
 NOR2_X1 _21596_ (.A1(_12011_),
    .A2(_11988_),
    .ZN(_12243_));
 OAI221_X1 _21597_ (.A(_14940_),
    .B1(_12008_),
    .B2(_12092_),
    .C1(_12243_),
    .C2(_12009_),
    .ZN(_12244_));
 NAND3_X1 _21598_ (.A1(net1014),
    .A2(_14922_),
    .A3(_12014_),
    .ZN(_12245_));
 NAND2_X1 _21599_ (.A1(_11914_),
    .A2(_11991_),
    .ZN(_12246_));
 OAI221_X1 _21600_ (.A(_14947_),
    .B1(_12050_),
    .B2(_12246_),
    .C1(_12041_),
    .C2(_14931_),
    .ZN(_12247_));
 NAND4_X1 _21601_ (.A1(_11998_),
    .A2(_12244_),
    .A3(_12245_),
    .A4(_12247_),
    .ZN(_12248_));
 NAND3_X1 _21602_ (.A1(_12004_),
    .A2(_12242_),
    .A3(_12248_),
    .ZN(_12249_));
 NOR2_X1 _21603_ (.A1(_11979_),
    .A2(_11974_),
    .ZN(_12250_));
 NAND2_X2 _21604_ (.A1(_11961_),
    .A2(_11912_),
    .ZN(_12251_));
 AOI21_X1 _21605_ (.A(_12251_),
    .B1(_11894_),
    .B2(_12153_),
    .ZN(_12252_));
 NAND2_X1 _21606_ (.A1(_11896_),
    .A2(_12017_),
    .ZN(_12253_));
 NOR2_X2 _21607_ (.A1(_12029_),
    .A2(_11895_),
    .ZN(_12254_));
 NOR2_X1 _21608_ (.A1(_12109_),
    .A2(_12254_),
    .ZN(_12255_));
 AOI21_X2 _21609_ (.A(_12098_),
    .B1(_12253_),
    .B2(_12255_),
    .ZN(_12256_));
 AOI221_X2 _21610_ (.A(_12003_),
    .B1(_12250_),
    .B2(_12252_),
    .C1(_12256_),
    .C2(_12231_),
    .ZN(_12257_));
 AOI21_X1 _21611_ (.A(_12023_),
    .B1(_12133_),
    .B2(_12118_),
    .ZN(_12258_));
 AOI21_X2 _21612_ (.A(_11990_),
    .B1(_12042_),
    .B2(_12176_),
    .ZN(_12259_));
 NOR3_X1 _21613_ (.A1(_12157_),
    .A2(_12258_),
    .A3(_12259_),
    .ZN(_12260_));
 OAI21_X1 _21614_ (.A(_14931_),
    .B1(_14947_),
    .B2(_12046_),
    .ZN(_12261_));
 AOI221_X2 _21615_ (.A(_12160_),
    .B1(_12010_),
    .B2(_11855_),
    .C1(_11916_),
    .C2(_12082_),
    .ZN(_12262_));
 AOI21_X1 _21616_ (.A(_12260_),
    .B1(_12261_),
    .B2(_12262_),
    .ZN(_12263_));
 AOI21_X1 _21617_ (.A(_11905_),
    .B1(_12257_),
    .B2(_12263_),
    .ZN(_12264_));
 NOR3_X2 _21618_ (.A1(_12052_),
    .A2(_12043_),
    .A3(_12136_),
    .ZN(_12265_));
 AOI221_X2 _21619_ (.A(_12265_),
    .B1(_12250_),
    .B2(net109),
    .C1(_12011_),
    .C2(_12082_),
    .ZN(_12266_));
 NAND2_X1 _21620_ (.A1(_12004_),
    .A2(_12266_),
    .ZN(_12267_));
 AOI21_X2 _21621_ (.A(_12163_),
    .B1(_12154_),
    .B2(_12084_),
    .ZN(_12268_));
 AOI21_X1 _21622_ (.A(net918),
    .B1(net1098),
    .B2(_12009_),
    .ZN(_12269_));
 AOI21_X1 _21623_ (.A(_12268_),
    .B1(_12269_),
    .B2(_14940_),
    .ZN(_12270_));
 AOI21_X1 _21624_ (.A(_12006_),
    .B1(_12075_),
    .B2(_12270_),
    .ZN(_12271_));
 AND3_X1 _21625_ (.A1(_12080_),
    .A2(net981),
    .A3(_12110_),
    .ZN(_12272_));
 NOR3_X1 _21626_ (.A1(_14947_),
    .A2(_12050_),
    .A3(net918),
    .ZN(_12273_));
 OAI21_X1 _21627_ (.A(_12004_),
    .B1(_12272_),
    .B2(_12273_),
    .ZN(_12274_));
 AOI221_X2 _21628_ (.A(_12003_),
    .B1(_12062_),
    .B2(_12029_),
    .C1(_11979_),
    .C2(_12109_),
    .ZN(_12275_));
 NOR2_X1 _21629_ (.A1(_11998_),
    .A2(_12275_),
    .ZN(_12276_));
 AOI22_X2 _21630_ (.A1(_12267_),
    .A2(_12271_),
    .B1(_12274_),
    .B2(_12276_),
    .ZN(_12277_));
 NOR3_X1 _21631_ (.A1(_12043_),
    .A2(_12115_),
    .A3(_12114_),
    .ZN(_12278_));
 MUX2_X1 _21632_ (.A(_11915_),
    .B(_11976_),
    .S(_12020_),
    .Z(_12279_));
 AOI21_X1 _21633_ (.A(_12278_),
    .B1(_12279_),
    .B2(_11896_),
    .ZN(_12280_));
 AOI21_X2 _21634_ (.A(_12127_),
    .B1(_12020_),
    .B2(_12016_),
    .ZN(_12281_));
 AOI22_X1 _21635_ (.A1(_11872_),
    .A2(_12061_),
    .B1(_11990_),
    .B2(_12281_),
    .ZN(_12282_));
 MUX2_X1 _21636_ (.A(_12280_),
    .B(_12282_),
    .S(_11962_),
    .Z(_12283_));
 NAND2_X1 _21637_ (.A1(_11976_),
    .A2(_11894_),
    .ZN(_12284_));
 NAND3_X1 _21638_ (.A1(_12021_),
    .A2(_11966_),
    .A3(_12284_),
    .ZN(_12285_));
 OAI21_X1 _21639_ (.A(_12074_),
    .B1(_12285_),
    .B2(_12006_),
    .ZN(_12286_));
 NOR2_X1 _21640_ (.A1(_11990_),
    .A2(_11961_),
    .ZN(_12287_));
 AOI22_X1 _21641_ (.A1(_12069_),
    .A2(_12101_),
    .B1(_12287_),
    .B2(_12021_),
    .ZN(_12288_));
 NOR2_X1 _21642_ (.A1(_12011_),
    .A2(_12288_),
    .ZN(_12289_));
 OAI33_X1 _21643_ (.A1(_12014_),
    .A2(_12075_),
    .A3(_12283_),
    .B1(_12286_),
    .B2(_12289_),
    .B3(_12036_),
    .ZN(_12290_));
 AOI222_X2 _21644_ (.A1(_12249_),
    .A2(_12264_),
    .B1(_12277_),
    .B2(_12060_),
    .C1(_12290_),
    .C2(_11905_),
    .ZN(_00067_));
 NOR2_X1 _21645_ (.A1(_12058_),
    .A2(_12003_),
    .ZN(_12291_));
 MUX2_X1 _21646_ (.A(_14936_),
    .B(_11971_),
    .S(_11968_),
    .Z(_12292_));
 OAI21_X1 _21647_ (.A(_12291_),
    .B1(_12292_),
    .B2(_12160_),
    .ZN(_12293_));
 INV_X1 _21648_ (.A(_12029_),
    .ZN(_12294_));
 OAI21_X4 _21649_ (.A(_11893_),
    .B1(_11943_),
    .B2(_11945_),
    .ZN(_12295_));
 AOI21_X1 _21650_ (.A(_12032_),
    .B1(_12019_),
    .B2(net2),
    .ZN(_12296_));
 OAI222_X2 _21651_ (.A1(_12294_),
    .A2(_12295_),
    .B1(_12084_),
    .B2(_12052_),
    .C1(_12296_),
    .C2(_11893_),
    .ZN(_12297_));
 NAND3_X1 _21652_ (.A1(_11915_),
    .A2(_11926_),
    .A3(_11931_),
    .ZN(_12298_));
 NAND2_X1 _21653_ (.A1(_12167_),
    .A2(_12298_),
    .ZN(_12299_));
 AOI221_X2 _21654_ (.A(_12239_),
    .B1(_12030_),
    .B2(_12061_),
    .C1(_12299_),
    .C2(_11989_),
    .ZN(_12300_));
 MUX2_X1 _21655_ (.A(_12297_),
    .B(_12300_),
    .S(_11987_),
    .Z(_12301_));
 AOI22_X2 _21656_ (.A1(_14928_),
    .A2(_12136_),
    .B1(_12176_),
    .B2(_12080_),
    .ZN(_12302_));
 AOI221_X2 _21657_ (.A(_12293_),
    .B1(_11963_),
    .B2(_12301_),
    .C1(_12158_),
    .C2(_12302_),
    .ZN(_12303_));
 OAI21_X1 _21658_ (.A(_11896_),
    .B1(_11975_),
    .B2(_12153_),
    .ZN(_12304_));
 AND2_X1 _21659_ (.A1(_12042_),
    .A2(_12176_),
    .ZN(_12305_));
 OAI221_X1 _21660_ (.A(_11988_),
    .B1(_12239_),
    .B2(_12304_),
    .C1(_12305_),
    .C2(_12023_),
    .ZN(_12306_));
 NAND2_X1 _21661_ (.A1(_12029_),
    .A2(_11895_),
    .ZN(_12307_));
 OAI21_X2 _21662_ (.A(_12307_),
    .B1(_12143_),
    .B2(_12023_),
    .ZN(_12308_));
 OAI21_X1 _21663_ (.A(_12306_),
    .B1(_12308_),
    .B2(_12008_),
    .ZN(_12309_));
 AND4_X2 _21664_ (.A1(_12309_),
    .A2(_11905_),
    .A3(_12004_),
    .A4(_12007_),
    .ZN(_12310_));
 NAND2_X1 _21665_ (.A1(net1144),
    .A2(_12136_),
    .ZN(_12311_));
 AOI21_X1 _21666_ (.A(_11989_),
    .B1(_11967_),
    .B2(_11915_),
    .ZN(_12312_));
 AOI21_X1 _21667_ (.A(_12142_),
    .B1(_11974_),
    .B2(net842),
    .ZN(_12313_));
 AOI221_X2 _21668_ (.A(_11913_),
    .B1(_12311_),
    .B2(_12312_),
    .C1(_12313_),
    .C2(_11990_),
    .ZN(_12314_));
 NAND2_X1 _21669_ (.A1(net1144),
    .A2(_12032_),
    .ZN(_12315_));
 NOR2_X1 _21670_ (.A1(_12069_),
    .A2(_12142_),
    .ZN(_12316_));
 MUX2_X1 _21671_ (.A(_12153_),
    .B(_12016_),
    .S(_11974_),
    .Z(_12317_));
 AOI22_X1 _21672_ (.A1(_12315_),
    .A2(_12316_),
    .B1(_12317_),
    .B2(_12080_),
    .ZN(_12318_));
 AOI21_X1 _21673_ (.A(_12314_),
    .B1(_12318_),
    .B2(_12041_),
    .ZN(_12319_));
 NOR4_X2 _21674_ (.A1(_12319_),
    .A2(_12059_),
    .A3(_12075_),
    .A4(_12007_),
    .ZN(_12320_));
 NAND2_X1 _21675_ (.A1(net978),
    .A2(_11965_),
    .ZN(_12321_));
 AOI21_X1 _21676_ (.A(_11975_),
    .B1(_12045_),
    .B2(_12321_),
    .ZN(_12322_));
 NOR3_X1 _21677_ (.A1(_11914_),
    .A2(_11984_),
    .A3(_12322_),
    .ZN(_12323_));
 NOR3_X1 _21678_ (.A1(_14940_),
    .A2(_11988_),
    .A3(_12121_),
    .ZN(_12324_));
 NOR3_X1 _21679_ (.A1(_12323_),
    .A2(_11998_),
    .A3(_12324_),
    .ZN(_12325_));
 NAND3_X1 _21680_ (.A1(_11916_),
    .A2(_11926_),
    .A3(_11931_),
    .ZN(_12326_));
 AND3_X1 _21681_ (.A1(_12163_),
    .A2(_11946_),
    .A3(_12326_),
    .ZN(_12327_));
 NOR3_X2 _21682_ (.A1(_12111_),
    .A2(_12251_),
    .A3(_12327_),
    .ZN(_12328_));
 NOR2_X1 _21683_ (.A1(_11904_),
    .A2(_12003_),
    .ZN(_12329_));
 OAI22_X1 _21684_ (.A1(_12153_),
    .A2(_11933_),
    .B1(_12136_),
    .B2(_12080_),
    .ZN(_12330_));
 OAI21_X1 _21685_ (.A(_12329_),
    .B1(_12330_),
    .B2(_12165_),
    .ZN(_12331_));
 AOI21_X2 _21686_ (.A(_11891_),
    .B1(_11967_),
    .B2(_11853_),
    .ZN(_12332_));
 AOI221_X2 _21687_ (.A(_11912_),
    .B1(_12298_),
    .B2(_12332_),
    .C1(_11965_),
    .C2(_14931_),
    .ZN(_12333_));
 NAND2_X2 _21688_ (.A1(_12030_),
    .A2(_12019_),
    .ZN(_12334_));
 AOI221_X1 _21689_ (.A(_11986_),
    .B1(_11974_),
    .B2(_12029_),
    .C1(_12334_),
    .C2(_12043_),
    .ZN(_12335_));
 NOR3_X1 _21690_ (.A1(_12335_),
    .A2(_12333_),
    .A3(_11963_),
    .ZN(_12336_));
 MUX2_X1 _21691_ (.A(_11893_),
    .B(_12133_),
    .S(_11986_),
    .Z(_12337_));
 NOR2_X1 _21692_ (.A1(_11855_),
    .A2(_12337_),
    .ZN(_12338_));
 NAND3_X1 _21693_ (.A1(_12016_),
    .A2(_11965_),
    .A3(_11987_),
    .ZN(_12339_));
 NAND2_X1 _21694_ (.A1(_11913_),
    .A2(_12105_),
    .ZN(_12340_));
 AOI21_X1 _21695_ (.A(_12109_),
    .B1(_12339_),
    .B2(_12340_),
    .ZN(_12341_));
 AOI21_X1 _21696_ (.A(_11874_),
    .B1(_11893_),
    .B2(_11986_),
    .ZN(_12342_));
 NOR3_X1 _21697_ (.A1(_11975_),
    .A2(_12044_),
    .A3(_12342_),
    .ZN(_12343_));
 NOR4_X1 _21698_ (.A1(_12006_),
    .A2(_12338_),
    .A3(_12341_),
    .A4(_12343_),
    .ZN(_12344_));
 NAND2_X1 _21699_ (.A1(_12059_),
    .A2(_12003_),
    .ZN(_12345_));
 OAI33_X1 _21700_ (.A1(_12325_),
    .A2(_12328_),
    .A3(_12331_),
    .B1(_12336_),
    .B2(_12344_),
    .B3(_12345_),
    .ZN(_12346_));
 NOR4_X4 _21701_ (.A1(_12346_),
    .A2(_12303_),
    .A3(_12320_),
    .A4(_12310_),
    .ZN(_00068_));
 OAI221_X2 _21702_ (.A(_12069_),
    .B1(_11975_),
    .B2(_12029_),
    .C1(_12133_),
    .C2(net715),
    .ZN(_12347_));
 AOI21_X1 _21703_ (.A(net1012),
    .B1(_12031_),
    .B2(net109),
    .ZN(_12348_));
 AOI21_X1 _21704_ (.A(_11903_),
    .B1(_12348_),
    .B2(_12163_),
    .ZN(_12349_));
 NOR2_X2 _21705_ (.A1(_11996_),
    .A2(_11965_),
    .ZN(_12350_));
 OAI22_X2 _21706_ (.A1(_12153_),
    .A2(_12295_),
    .B1(_12350_),
    .B2(_12009_),
    .ZN(_12351_));
 AOI221_X2 _21707_ (.A(_12008_),
    .B1(_12349_),
    .B2(_12347_),
    .C1(_12351_),
    .C2(_11904_),
    .ZN(_12352_));
 OAI21_X1 _21708_ (.A(net1014),
    .B1(_14922_),
    .B2(_12061_),
    .ZN(_12353_));
 AOI21_X1 _21709_ (.A(_11905_),
    .B1(_12133_),
    .B2(_12353_),
    .ZN(_12354_));
 AOI21_X1 _21710_ (.A(_11979_),
    .B1(_11983_),
    .B2(_11903_),
    .ZN(_12355_));
 NAND2_X1 _21711_ (.A1(_11967_),
    .A2(_11902_),
    .ZN(_12356_));
 OAI221_X1 _21712_ (.A(_12014_),
    .B1(_12110_),
    .B2(_12355_),
    .C1(_12356_),
    .C2(_12253_),
    .ZN(_12357_));
 OAI21_X1 _21713_ (.A(_12075_),
    .B1(_12354_),
    .B2(_12357_),
    .ZN(_12358_));
 INV_X1 _21714_ (.A(_12254_),
    .ZN(_12359_));
 AOI21_X1 _21715_ (.A(_11968_),
    .B1(_12015_),
    .B2(_12016_),
    .ZN(_12360_));
 AOI21_X2 _21716_ (.A(_12036_),
    .B1(_12359_),
    .B2(_12360_),
    .ZN(_12361_));
 AOI21_X1 _21717_ (.A(_11894_),
    .B1(_11936_),
    .B2(_11946_),
    .ZN(_12362_));
 NOR2_X1 _21718_ (.A1(_11914_),
    .A2(_12362_),
    .ZN(_12363_));
 AOI221_X2 _21719_ (.A(_11904_),
    .B1(_12361_),
    .B2(_11946_),
    .C1(_12363_),
    .C2(_12081_),
    .ZN(_12364_));
 OAI22_X1 _21720_ (.A1(_12120_),
    .A2(_12009_),
    .B1(_12010_),
    .B2(_14928_),
    .ZN(_12365_));
 OAI221_X2 _21721_ (.A(_12076_),
    .B1(_12214_),
    .B2(_14931_),
    .C1(_12064_),
    .C2(_12295_),
    .ZN(_12366_));
 NAND2_X1 _21722_ (.A1(_14928_),
    .A2(_12082_),
    .ZN(_12367_));
 AOI21_X1 _21723_ (.A(_14922_),
    .B1(_12053_),
    .B2(_12367_),
    .ZN(_12368_));
 OAI221_X2 _21724_ (.A(_12004_),
    .B1(_12100_),
    .B2(_12365_),
    .C1(_12366_),
    .C2(_12368_),
    .ZN(_12369_));
 OAI22_X2 _21725_ (.A1(_12352_),
    .A2(_12358_),
    .B1(_12369_),
    .B2(_12364_),
    .ZN(_12370_));
 NOR2_X1 _21726_ (.A1(_11965_),
    .A2(_12167_),
    .ZN(_12371_));
 AND2_X1 _21727_ (.A1(_12163_),
    .A2(_12305_),
    .ZN(_12372_));
 OAI21_X1 _21728_ (.A(_12059_),
    .B1(_12371_),
    .B2(_12372_),
    .ZN(_12373_));
 NOR2_X1 _21729_ (.A1(net1199),
    .A2(_12035_),
    .ZN(_12374_));
 OAI21_X1 _21730_ (.A(_12118_),
    .B1(_12031_),
    .B2(_11915_),
    .ZN(_12375_));
 AOI21_X1 _21731_ (.A(_12374_),
    .B1(_12375_),
    .B2(_12069_),
    .ZN(_12376_));
 AOI21_X1 _21732_ (.A(_11914_),
    .B1(_11904_),
    .B2(_12376_),
    .ZN(_12377_));
 AOI221_X2 _21733_ (.A(_11902_),
    .B1(_12315_),
    .B2(_11893_),
    .C1(_12031_),
    .C2(net978),
    .ZN(_12378_));
 NOR2_X1 _21734_ (.A1(_12014_),
    .A2(_12378_),
    .ZN(_12379_));
 AND2_X1 _21735_ (.A1(_11992_),
    .A2(_11936_),
    .ZN(_12380_));
 OAI221_X2 _21736_ (.A(_11904_),
    .B1(_12214_),
    .B2(_14928_),
    .C1(_12380_),
    .C2(_14940_),
    .ZN(_12381_));
 AOI221_X2 _21737_ (.A(_12075_),
    .B1(_12373_),
    .B2(_12377_),
    .C1(_12379_),
    .C2(_12381_),
    .ZN(_12382_));
 OAI221_X2 _21738_ (.A(_12060_),
    .B1(_12214_),
    .B2(_12120_),
    .C1(_12022_),
    .C2(_12064_),
    .ZN(_12383_));
 NOR3_X4 _21739_ (.A1(_11943_),
    .A2(_11970_),
    .A3(_11945_),
    .ZN(_12384_));
 NOR3_X2 _21740_ (.A1(_14947_),
    .A2(_12384_),
    .A3(net1012),
    .ZN(_12385_));
 OAI21_X1 _21741_ (.A(_12118_),
    .B1(_12031_),
    .B2(_11976_),
    .ZN(_12386_));
 AOI21_X2 _21742_ (.A(_12385_),
    .B1(_12386_),
    .B2(_14947_),
    .ZN(_12387_));
 OAI211_X2 _21743_ (.A(_12075_),
    .B(_12383_),
    .C1(_12095_),
    .C2(_12387_),
    .ZN(_12388_));
 OAI21_X1 _21744_ (.A(_12021_),
    .B1(_12350_),
    .B2(_11979_),
    .ZN(_12389_));
 AOI22_X1 _21745_ (.A1(_12120_),
    .A2(_12061_),
    .B1(_12386_),
    .B2(_12069_),
    .ZN(_12390_));
 AOI221_X2 _21746_ (.A(_11904_),
    .B1(_12389_),
    .B2(_11995_),
    .C1(_12390_),
    .C2(_11914_),
    .ZN(_12391_));
 OAI21_X2 _21747_ (.A(_11998_),
    .B1(_12388_),
    .B2(_12391_),
    .ZN(_12392_));
 OAI22_X2 _21748_ (.A1(_12370_),
    .A2(_11998_),
    .B1(_12382_),
    .B2(_12392_),
    .ZN(_00069_));
 NOR2_X1 _21749_ (.A1(_12153_),
    .A2(_11894_),
    .ZN(_12393_));
 AOI22_X1 _21750_ (.A1(_11988_),
    .A2(_12025_),
    .B1(_12393_),
    .B2(_12021_),
    .ZN(_12394_));
 NAND2_X1 _21751_ (.A1(_11874_),
    .A2(_12043_),
    .ZN(_12395_));
 NAND2_X1 _21752_ (.A1(_12008_),
    .A2(_12009_),
    .ZN(_12396_));
 OAI221_X1 _21753_ (.A(_12329_),
    .B1(_12394_),
    .B2(net1014),
    .C1(_12395_),
    .C2(_12396_),
    .ZN(_12397_));
 AOI21_X1 _21754_ (.A(_12115_),
    .B1(_12015_),
    .B2(net1014),
    .ZN(_12398_));
 OAI221_X1 _21755_ (.A(_12025_),
    .B1(_12133_),
    .B2(_14928_),
    .C1(_12398_),
    .C2(_12153_),
    .ZN(_12399_));
 AOI22_X1 _21756_ (.A1(_12007_),
    .A2(_12397_),
    .B1(_12399_),
    .B2(_12140_),
    .ZN(_12400_));
 OAI21_X1 _21757_ (.A(_12041_),
    .B1(_12374_),
    .B2(_12268_),
    .ZN(_12401_));
 MUX2_X1 _21758_ (.A(_12294_),
    .B(net1013),
    .S(_12163_),
    .Z(_12402_));
 MUX2_X1 _21759_ (.A(_14942_),
    .B(_12402_),
    .S(_12022_),
    .Z(_12403_));
 OAI21_X2 _21760_ (.A(_12401_),
    .B1(_12403_),
    .B2(_12041_),
    .ZN(_12404_));
 AOI21_X1 _21761_ (.A(_12400_),
    .B1(_12404_),
    .B2(_12291_),
    .ZN(_12405_));
 NOR2_X1 _21762_ (.A1(_11968_),
    .A2(_12058_),
    .ZN(_12406_));
 MUX2_X1 _21763_ (.A(_11969_),
    .B(_14932_),
    .S(_11912_),
    .Z(_12407_));
 OR2_X1 _21764_ (.A1(_11893_),
    .A2(_12017_),
    .ZN(_12408_));
 OAI221_X1 _21765_ (.A(_12406_),
    .B1(_12407_),
    .B2(_11965_),
    .C1(_12408_),
    .C2(_11913_),
    .ZN(_12409_));
 AOI21_X1 _21766_ (.A(net1144),
    .B1(_11874_),
    .B2(_11986_),
    .ZN(_12410_));
 NAND2_X1 _21767_ (.A1(_11872_),
    .A2(_11892_),
    .ZN(_12411_));
 NOR2_X1 _21768_ (.A1(_11912_),
    .A2(_12411_),
    .ZN(_12412_));
 OR4_X1 _21769_ (.A1(_11979_),
    .A2(_12356_),
    .A3(_12410_),
    .A4(_12412_),
    .ZN(_12413_));
 AND3_X1 _21770_ (.A1(_12003_),
    .A2(_12409_),
    .A3(_12413_),
    .ZN(_12414_));
 AND2_X1 _21771_ (.A1(_11892_),
    .A2(_11991_),
    .ZN(_12415_));
 NAND2_X1 _21772_ (.A1(_14926_),
    .A2(_11967_),
    .ZN(_12416_));
 AND2_X1 _21773_ (.A1(_11891_),
    .A2(_12118_),
    .ZN(_12417_));
 AOI221_X2 _21774_ (.A(_11912_),
    .B1(_12161_),
    .B2(_12415_),
    .C1(_12416_),
    .C2(_12417_),
    .ZN(_12418_));
 NAND2_X2 _21775_ (.A1(_11989_),
    .A2(_12017_),
    .ZN(_12419_));
 OAI221_X2 _21776_ (.A(_11912_),
    .B1(_12419_),
    .B2(_12019_),
    .C1(_11932_),
    .C2(_11970_),
    .ZN(_12420_));
 OAI21_X1 _21777_ (.A(_12084_),
    .B1(_12020_),
    .B2(_12029_),
    .ZN(_12421_));
 AOI21_X2 _21778_ (.A(_12420_),
    .B1(_12421_),
    .B2(_12043_),
    .ZN(_12422_));
 OR3_X4 _21779_ (.A1(_12422_),
    .A2(_12418_),
    .A3(_11903_),
    .ZN(_12423_));
 MUX2_X1 _21780_ (.A(_12029_),
    .B(_12064_),
    .S(_12020_),
    .Z(_12424_));
 OAI221_X1 _21781_ (.A(_12076_),
    .B1(_12424_),
    .B2(_12023_),
    .C1(_12065_),
    .C2(_14928_),
    .ZN(_12425_));
 OAI21_X1 _21782_ (.A(_12058_),
    .B1(_12295_),
    .B2(_14931_),
    .ZN(_12426_));
 OAI221_X2 _21783_ (.A(_11988_),
    .B1(_12149_),
    .B2(_12356_),
    .C1(_12426_),
    .C2(_12259_),
    .ZN(_12427_));
 OAI21_X1 _21784_ (.A(_12065_),
    .B1(_12163_),
    .B2(_11855_),
    .ZN(_12428_));
 OAI21_X1 _21785_ (.A(_12085_),
    .B1(_12428_),
    .B2(_12115_),
    .ZN(_12429_));
 NAND3_X2 _21786_ (.A1(_12429_),
    .A2(_12427_),
    .A3(_12425_),
    .ZN(_12430_));
 AOI221_X2 _21787_ (.A(_12007_),
    .B1(_12423_),
    .B2(_12414_),
    .C1(_12430_),
    .C2(_12075_),
    .ZN(_12431_));
 OAI21_X1 _21788_ (.A(_11904_),
    .B1(_12022_),
    .B2(_14943_),
    .ZN(_12432_));
 MUX2_X1 _21789_ (.A(_12011_),
    .B(_12229_),
    .S(_12080_),
    .Z(_12433_));
 AOI21_X1 _21790_ (.A(_12432_),
    .B1(_12433_),
    .B2(_12022_),
    .ZN(_12434_));
 NAND2_X1 _21791_ (.A1(_12326_),
    .A2(_12176_),
    .ZN(_12435_));
 AOI221_X2 _21792_ (.A(_11903_),
    .B1(_12435_),
    .B2(_12163_),
    .C1(_11982_),
    .C2(_14926_),
    .ZN(_12436_));
 NOR3_X1 _21793_ (.A1(_12014_),
    .A2(_12434_),
    .A3(_12436_),
    .ZN(_12437_));
 NOR2_X1 _21794_ (.A1(_12161_),
    .A2(_12194_),
    .ZN(_12438_));
 OR3_X1 _21795_ (.A1(_14941_),
    .A2(_14950_),
    .A3(_11975_),
    .ZN(_12439_));
 NAND3_X1 _21796_ (.A1(_12014_),
    .A2(_12059_),
    .A3(_12439_),
    .ZN(_12440_));
 AOI211_X2 _21797_ (.A(_11990_),
    .B(_12384_),
    .C1(_11975_),
    .C2(net109),
    .ZN(_12441_));
 AOI21_X1 _21798_ (.A(_12441_),
    .B1(_12033_),
    .B2(_14947_),
    .ZN(_12442_));
 OAI22_X1 _21799_ (.A1(_12438_),
    .A2(_12440_),
    .B1(_12442_),
    .B2(_12100_),
    .ZN(_12443_));
 OAI21_X1 _21800_ (.A(_12004_),
    .B1(_12437_),
    .B2(_12443_),
    .ZN(_12444_));
 AOI21_X1 _21801_ (.A(_12007_),
    .B1(_12414_),
    .B2(_12423_),
    .ZN(_12445_));
 OAI22_X1 _21802_ (.A1(_12431_),
    .A2(_12405_),
    .B1(_12444_),
    .B2(_12445_),
    .ZN(_00070_));
 AOI211_X2 _21803_ (.A(_11989_),
    .B(_12114_),
    .C1(_12019_),
    .C2(net1144),
    .ZN(_12446_));
 OAI21_X2 _21804_ (.A(_11964_),
    .B1(_12128_),
    .B2(_12446_),
    .ZN(_12447_));
 NOR2_X1 _21805_ (.A1(_14950_),
    .A2(_12031_),
    .ZN(_12448_));
 AND3_X1 _21806_ (.A1(_12020_),
    .A2(_12045_),
    .A3(_12307_),
    .ZN(_12449_));
 OAI21_X1 _21807_ (.A(_11987_),
    .B1(_12448_),
    .B2(_12449_),
    .ZN(_12450_));
 AND3_X4 _21808_ (.A1(_12447_),
    .A2(_11962_),
    .A3(_12450_),
    .ZN(_12451_));
 NOR2_X1 _21809_ (.A1(_14936_),
    .A2(_12109_),
    .ZN(_12452_));
 NOR3_X1 _21810_ (.A1(_12030_),
    .A2(_11965_),
    .A3(_11968_),
    .ZN(_12453_));
 OAI21_X1 _21811_ (.A(_11988_),
    .B1(_12452_),
    .B2(_12453_),
    .ZN(_12454_));
 MUX2_X1 _21812_ (.A(_11937_),
    .B(_11853_),
    .S(_11989_),
    .Z(_12455_));
 NAND2_X1 _21813_ (.A1(_12395_),
    .A2(_12031_),
    .ZN(_12456_));
 OAI221_X2 _21814_ (.A(_11964_),
    .B1(_12109_),
    .B2(_12455_),
    .C1(_12456_),
    .C2(net1013),
    .ZN(_12457_));
 AOI21_X2 _21815_ (.A(_11963_),
    .B1(_12454_),
    .B2(_12457_),
    .ZN(_12458_));
 NOR4_X4 _21816_ (.A1(_12458_),
    .A2(_12075_),
    .A3(_12451_),
    .A4(_12059_),
    .ZN(_12459_));
 NAND2_X1 _21817_ (.A1(_11904_),
    .A2(_12074_),
    .ZN(_12460_));
 MUX2_X1 _21818_ (.A(_12010_),
    .B(_12082_),
    .S(_11872_),
    .Z(_12461_));
 AOI221_X2 _21819_ (.A(_12251_),
    .B1(_12461_),
    .B2(_11855_),
    .C1(_12061_),
    .C2(net1199),
    .ZN(_12462_));
 NOR2_X1 _21820_ (.A1(_12120_),
    .A2(_12109_),
    .ZN(_12463_));
 NOR4_X1 _21821_ (.A1(_14947_),
    .A2(_12384_),
    .A3(_12463_),
    .A4(_12165_),
    .ZN(_12464_));
 NOR3_X1 _21822_ (.A1(_12460_),
    .A2(_12462_),
    .A3(_12464_),
    .ZN(_12465_));
 NAND2_X1 _21823_ (.A1(_11933_),
    .A2(_12167_),
    .ZN(_12466_));
 NAND2_X1 _21824_ (.A1(net1013),
    .A2(_12466_),
    .ZN(_12467_));
 AOI21_X1 _21825_ (.A(_11914_),
    .B1(_12311_),
    .B2(_12467_),
    .ZN(_12468_));
 AOI21_X1 _21826_ (.A(_11982_),
    .B1(_12021_),
    .B2(_11979_),
    .ZN(_12469_));
 AOI21_X1 _21827_ (.A(_12115_),
    .B1(_12082_),
    .B2(_14922_),
    .ZN(_12470_));
 OAI22_X1 _21828_ (.A1(net1014),
    .A2(_12469_),
    .B1(_12470_),
    .B2(_11988_),
    .ZN(_12471_));
 OAI21_X1 _21829_ (.A(_12007_),
    .B1(_12468_),
    .B2(_12471_),
    .ZN(_12472_));
 NAND2_X1 _21830_ (.A1(net1144),
    .A2(_11974_),
    .ZN(_12473_));
 AOI221_X2 _21831_ (.A(_11964_),
    .B1(_12473_),
    .B2(_12415_),
    .C1(_12213_),
    .C2(_12023_),
    .ZN(_12474_));
 OAI222_X2 _21832_ (.A1(_14931_),
    .A2(_11933_),
    .B1(_12065_),
    .B2(_12153_),
    .C1(_12011_),
    .C2(_12062_),
    .ZN(_12475_));
 NOR2_X1 _21833_ (.A1(_12014_),
    .A2(_12475_),
    .ZN(_12476_));
 OAI21_X1 _21834_ (.A(_12057_),
    .B1(_12474_),
    .B2(_12476_),
    .ZN(_12477_));
 AOI221_X2 _21835_ (.A(_12005_),
    .B1(_12334_),
    .B2(_12332_),
    .C1(_11895_),
    .C2(_11916_),
    .ZN(_12478_));
 AOI22_X1 _21836_ (.A1(_11976_),
    .A2(_11974_),
    .B1(_12115_),
    .B2(_11853_),
    .ZN(_12479_));
 NOR3_X1 _21837_ (.A1(_11896_),
    .A2(_11961_),
    .A3(_12479_),
    .ZN(_12480_));
 NOR2_X1 _21838_ (.A1(_11913_),
    .A2(_12074_),
    .ZN(_12481_));
 OAI21_X1 _21839_ (.A(_12481_),
    .B1(_12171_),
    .B2(_11962_),
    .ZN(_12482_));
 OR3_X1 _21840_ (.A1(_12478_),
    .A2(_12480_),
    .A3(_12482_),
    .ZN(_12483_));
 OR2_X1 _21841_ (.A1(_12161_),
    .A2(_12194_),
    .ZN(_12484_));
 NOR3_X2 _21842_ (.A1(_12142_),
    .A2(_12074_),
    .A3(_12251_),
    .ZN(_12485_));
 NAND2_X1 _21843_ (.A1(_12473_),
    .A2(_12417_),
    .ZN(_12486_));
 NAND3_X1 _21844_ (.A1(_12005_),
    .A2(_11986_),
    .A3(_12074_),
    .ZN(_12487_));
 AOI21_X1 _21845_ (.A(_12487_),
    .B1(_12254_),
    .B2(_11974_),
    .ZN(_12488_));
 AOI221_X2 _21846_ (.A(_11903_),
    .B1(_12485_),
    .B2(_12484_),
    .C1(_12486_),
    .C2(_12488_),
    .ZN(_12489_));
 OAI21_X1 _21847_ (.A(_11855_),
    .B1(_12136_),
    .B2(_12371_),
    .ZN(_12490_));
 AOI22_X1 _21848_ (.A1(_11872_),
    .A2(_12010_),
    .B1(_12082_),
    .B2(_11915_),
    .ZN(_12491_));
 NAND4_X1 _21849_ (.A1(_12074_),
    .A2(_12140_),
    .A3(_12490_),
    .A4(_12491_),
    .ZN(_12492_));
 OAI221_X1 _21850_ (.A(_12053_),
    .B1(_12421_),
    .B2(_11896_),
    .C1(net1100),
    .C2(_12065_),
    .ZN(_12493_));
 NAND3_X1 _21851_ (.A1(_12003_),
    .A2(_12140_),
    .A3(_12493_),
    .ZN(_12494_));
 AND4_X2 _21852_ (.A1(_12489_),
    .A2(_12483_),
    .A3(_12492_),
    .A4(_12494_),
    .ZN(_12495_));
 AOI221_X2 _21853_ (.A(_12459_),
    .B1(_12465_),
    .B2(_12472_),
    .C1(_12477_),
    .C2(_12495_),
    .ZN(_00071_));
 NAND2_X1 _21854_ (.A1(_06256_),
    .A2(_09023_),
    .ZN(_12496_));
 OR2_X1 _21855_ (.A1(_06256_),
    .A2(_09015_),
    .ZN(_12497_));
 XNOR2_X2 _21856_ (.A(\sa01_sr[1] ),
    .B(\sa30_sub[1] ),
    .ZN(_12498_));
 XNOR2_X2 _21857_ (.A(_09797_),
    .B(_12498_),
    .ZN(_12499_));
 XNOR2_X1 _21858_ (.A(_09739_),
    .B(net635),
    .ZN(_12500_));
 XNOR2_X1 _21859_ (.A(_12500_),
    .B(_12499_),
    .ZN(_12501_));
 MUX2_X2 _21860_ (.A(_12496_),
    .B(_12497_),
    .S(_12501_),
    .Z(_12502_));
 NOR3_X2 _21861_ (.A1(_06256_),
    .A2(_09194_),
    .A3(_00455_),
    .ZN(_12503_));
 AND2_X1 _21862_ (.A1(_06256_),
    .A2(_09727_),
    .ZN(_12504_));
 AOI21_X4 _21863_ (.A(_12503_),
    .B1(_12504_),
    .B2(_00455_),
    .ZN(_12505_));
 AND2_X4 _21864_ (.A1(_12502_),
    .A2(_12505_),
    .ZN(_12506_));
 BUF_X4 clone139 (.A(_12506_),
    .Z(net139));
 INV_X8 _21866_ (.A(_12506_),
    .ZN(_12508_));
 BUF_X1 rebuffer563 (.A(_06368_),
    .Z(net1162));
 BUF_X32 _21868_ (.A(_12508_),
    .Z(_14960_));
 XNOR2_X2 _21869_ (.A(_09719_),
    .B(\sa30_sub[0] ),
    .ZN(_12510_));
 XNOR2_X1 _21870_ (.A(net760),
    .B(_12510_),
    .ZN(_12511_));
 XOR2_X2 _21871_ (.A(net616),
    .B(_09796_),
    .Z(_12512_));
 NAND3_X1 _21872_ (.A1(_06242_),
    .A2(_09012_),
    .A3(_12512_),
    .ZN(_12513_));
 NOR2_X1 _21873_ (.A1(_06242_),
    .A2(_09015_),
    .ZN(_12514_));
 NAND2_X1 _21874_ (.A1(net670),
    .A2(_12514_),
    .ZN(_12515_));
 AOI21_X2 _21875_ (.A(_12511_),
    .B1(_12513_),
    .B2(_12515_),
    .ZN(_12516_));
 XOR2_X2 _21876_ (.A(\sa30_sub[0] ),
    .B(_09719_),
    .Z(_12517_));
 XNOR2_X1 _21877_ (.A(net760),
    .B(_12517_),
    .ZN(_12518_));
 NAND2_X1 _21878_ (.A1(_12512_),
    .A2(_12514_),
    .ZN(_12519_));
 NAND3_X1 _21879_ (.A1(_06242_),
    .A2(_09023_),
    .A3(net670),
    .ZN(_12520_));
 AOI21_X1 _21880_ (.A(_12518_),
    .B1(_12519_),
    .B2(_12520_),
    .ZN(_12521_));
 INV_X1 _21881_ (.A(_06242_),
    .ZN(_12522_));
 NAND3_X1 _21882_ (.A1(_12522_),
    .A2(_09028_),
    .A3(_00456_),
    .ZN(_12523_));
 NAND2_X1 _21883_ (.A1(_06242_),
    .A2(_09030_),
    .ZN(_12524_));
 OAI21_X1 _21884_ (.A(_12523_),
    .B1(_12524_),
    .B2(_00456_),
    .ZN(_12525_));
 OR3_X4 _21885_ (.A1(_12521_),
    .A2(_12516_),
    .A3(_12525_),
    .ZN(_12526_));
 INV_X8 _21886_ (.A(net606),
    .ZN(_12527_));
 BUF_X8 clone98 (.A(_06352_),
    .Z(net98));
 BUF_X8 _21888_ (.A(_12527_),
    .Z(_14963_));
 XNOR2_X2 _21889_ (.A(_09759_),
    .B(_09835_),
    .ZN(_12529_));
 XNOR2_X1 _21890_ (.A(_09763_),
    .B(_12529_),
    .ZN(_12530_));
 INV_X1 _21891_ (.A(_06297_),
    .ZN(_12531_));
 OR3_X1 _21892_ (.A1(_12531_),
    .A2(_08972_),
    .A3(net637),
    .ZN(_12532_));
 NAND3_X1 _21893_ (.A1(_12531_),
    .A2(_09099_),
    .A3(net638),
    .ZN(_12533_));
 AOI21_X2 _21894_ (.A(_12530_),
    .B1(_12532_),
    .B2(_12533_),
    .ZN(_12534_));
 XOR2_X2 _21895_ (.A(_09759_),
    .B(_09835_),
    .Z(_12535_));
 XNOR2_X1 _21896_ (.A(_09763_),
    .B(_12535_),
    .ZN(_12536_));
 OR3_X1 _21897_ (.A1(_06297_),
    .A2(_08992_),
    .A3(net637),
    .ZN(_12537_));
 NAND3_X1 _21898_ (.A1(_06297_),
    .A2(net947),
    .A3(net637),
    .ZN(_12538_));
 AOI21_X2 _21899_ (.A(_12536_),
    .B1(_12537_),
    .B2(_12538_),
    .ZN(_12539_));
 NAND3_X1 _21900_ (.A1(_12531_),
    .A2(_09015_),
    .A3(_00457_),
    .ZN(_12540_));
 NAND2_X1 _21901_ (.A1(_06297_),
    .A2(_09015_),
    .ZN(_12541_));
 OAI21_X2 _21902_ (.A(_12540_),
    .B1(_12541_),
    .B2(_00457_),
    .ZN(_12542_));
 NOR3_X4 _21903_ (.A1(_12534_),
    .A2(_12539_),
    .A3(_12542_),
    .ZN(_12543_));
 INV_X4 _21904_ (.A(_12543_),
    .ZN(_12544_));
 BUF_X4 _21905_ (.A(_12544_),
    .Z(_12545_));
 BUF_X4 _21906_ (.A(_12545_),
    .Z(_12546_));
 BUF_X4 _21907_ (.A(_12546_),
    .Z(_12547_));
 BUF_X4 _21908_ (.A(_12547_),
    .Z(_14979_));
 BUF_X16 _21909_ (.A(_12526_),
    .Z(_12548_));
 BUF_X8 _21910_ (.A(_12548_),
    .Z(_12549_));
 BUF_X8 _21911_ (.A(_12549_),
    .Z(_14954_));
 BUF_X4 _21912_ (.A(_12543_),
    .Z(_12550_));
 BUF_X4 _21913_ (.A(_12550_),
    .Z(_12551_));
 BUF_X4 _21914_ (.A(_12551_),
    .Z(_12552_));
 BUF_X4 _21915_ (.A(_12552_),
    .Z(_14972_));
 INV_X1 _21916_ (.A(_06282_),
    .ZN(_12553_));
 NOR2_X1 _21917_ (.A1(_12553_),
    .A2(_09028_),
    .ZN(_12554_));
 NOR2_X1 _21918_ (.A1(_06282_),
    .A2(_09028_),
    .ZN(_12555_));
 XNOR2_X1 _21919_ (.A(_09872_),
    .B(_09796_),
    .ZN(_12556_));
 XNOR2_X2 _21920_ (.A(_09836_),
    .B(_12556_),
    .ZN(_12557_));
 XOR2_X1 _21921_ (.A(_09869_),
    .B(_09813_),
    .Z(_12558_));
 XNOR2_X1 _21922_ (.A(_09840_),
    .B(_12558_),
    .ZN(_12559_));
 XNOR2_X1 _21923_ (.A(_12557_),
    .B(_12559_),
    .ZN(_12560_));
 MUX2_X2 _21924_ (.A(_12554_),
    .B(_12555_),
    .S(_12560_),
    .Z(_12561_));
 NAND3_X1 _21925_ (.A1(_12553_),
    .A2(_11938_),
    .A3(\text_in_r[84] ),
    .ZN(_12562_));
 NAND2_X1 _21926_ (.A1(_06282_),
    .A2(_11841_),
    .ZN(_12563_));
 OAI21_X4 _21927_ (.A(_12562_),
    .B1(_12563_),
    .B2(\text_in_r[84] ),
    .ZN(_12564_));
 OR2_X1 _21928_ (.A1(_12561_),
    .A2(_12564_),
    .ZN(_12565_));
 BUF_X4 _21929_ (.A(_12565_),
    .Z(_12566_));
 BUF_X4 _21930_ (.A(_12566_),
    .Z(_12567_));
 BUF_X4 _21931_ (.A(_12567_),
    .Z(_12568_));
 NAND2_X1 _21932_ (.A1(_08992_),
    .A2(\text_in_r[83] ),
    .ZN(_12569_));
 NAND3_X2 _21933_ (.A1(_06222_),
    .A2(_08974_),
    .A3(_12569_),
    .ZN(_12570_));
 OR2_X1 _21934_ (.A1(_06222_),
    .A2(_12569_),
    .ZN(_12571_));
 AND2_X2 _21935_ (.A1(_12570_),
    .A2(_12571_),
    .ZN(_12572_));
 NAND2_X1 _21936_ (.A1(_06222_),
    .A2(_12569_),
    .ZN(_12573_));
 OR2_X1 _21937_ (.A1(_06222_),
    .A2(_09727_),
    .ZN(_12574_));
 XNOR2_X2 _21938_ (.A(_09841_),
    .B(_09796_),
    .ZN(_12575_));
 XNOR2_X1 _21939_ (.A(_09764_),
    .B(_12575_),
    .ZN(_12576_));
 XOR2_X2 _21940_ (.A(_09836_),
    .B(_09868_),
    .Z(_12577_));
 XNOR2_X2 _21941_ (.A(net705),
    .B(_12577_),
    .ZN(_12578_));
 XNOR2_X2 _21942_ (.A(_12576_),
    .B(_12578_),
    .ZN(_12579_));
 MUX2_X2 _21943_ (.A(_12573_),
    .B(_12574_),
    .S(_12579_),
    .Z(_12580_));
 NAND2_X4 _21944_ (.A1(_12572_),
    .A2(_12580_),
    .ZN(_12581_));
 BUF_X4 _21945_ (.A(_12581_),
    .Z(_12582_));
 NOR2_X2 _21946_ (.A1(net723),
    .A2(_12582_),
    .ZN(_12583_));
 NAND2_X1 _21947_ (.A1(_14954_),
    .A2(_12547_),
    .ZN(_12584_));
 BUF_X4 clone146 (.A(net773),
    .Z(net146));
 NAND2_X4 _21949_ (.A1(_12570_),
    .A2(_12571_),
    .ZN(_12586_));
 AND2_X1 _21950_ (.A1(_06222_),
    .A2(_12569_),
    .ZN(_12587_));
 NOR2_X1 _21951_ (.A1(_06222_),
    .A2(_08973_),
    .ZN(_12588_));
 MUX2_X1 _21952_ (.A(_12587_),
    .B(_12588_),
    .S(_12579_),
    .Z(_12589_));
 BUF_X8 _21953_ (.A(_12589_),
    .Z(_12590_));
 NOR2_X4 _21954_ (.A1(_12586_),
    .A2(_12590_),
    .ZN(_12591_));
 BUF_X4 _21955_ (.A(_12591_),
    .Z(_12592_));
 BUF_X4 _21956_ (.A(_12592_),
    .Z(_12593_));
 MUX2_X1 _21957_ (.A(net138),
    .B(_14960_),
    .S(_12593_),
    .Z(_12594_));
 OAI221_X1 _21958_ (.A(_12568_),
    .B1(_12583_),
    .B2(_12584_),
    .C1(_12594_),
    .C2(_14979_),
    .ZN(_12595_));
 BUF_X8 _21959_ (.A(_12572_),
    .Z(_12596_));
 BUF_X8 _21960_ (.A(_12580_),
    .Z(_12597_));
 AOI21_X2 _21961_ (.A(_12543_),
    .B1(_12596_),
    .B2(_12597_),
    .ZN(_12598_));
 BUF_X4 _21962_ (.A(_12598_),
    .Z(_12599_));
 NAND2_X2 _21963_ (.A1(_12548_),
    .A2(_12599_),
    .ZN(_12600_));
 BUF_X4 _21964_ (.A(_12550_),
    .Z(_12601_));
 BUF_X4 _21965_ (.A(_12596_),
    .Z(_12602_));
 BUF_X8 _21966_ (.A(_12597_),
    .Z(_12603_));
 NAND3_X2 _21967_ (.A1(_12601_),
    .A2(_12602_),
    .A3(_12603_),
    .ZN(_12604_));
 BUF_X4 _21968_ (.A(_14958_),
    .Z(_12605_));
 BUF_X16 _21969_ (.A(_12506_),
    .Z(_12606_));
 BUF_X16 _21970_ (.A(_12606_),
    .Z(_14955_));
 NOR3_X4 _21971_ (.A1(_12550_),
    .A2(_12586_),
    .A3(_12590_),
    .ZN(_12607_));
 AOI21_X4 _21972_ (.A(_12544_),
    .B1(_12596_),
    .B2(_12597_),
    .ZN(_12608_));
 BUF_X4 _21973_ (.A(_12608_),
    .Z(_12609_));
 AOI21_X1 _21974_ (.A(_12607_),
    .B1(_12609_),
    .B2(_14963_),
    .ZN(_12610_));
 OAI221_X1 _21975_ (.A(_12600_),
    .B1(_12604_),
    .B2(_12605_),
    .C1(net200),
    .C2(_12610_),
    .ZN(_12611_));
 BUF_X4 _21976_ (.A(_12568_),
    .Z(_12612_));
 OAI21_X1 _21977_ (.A(_12595_),
    .B1(_12611_),
    .B2(_12612_),
    .ZN(_12613_));
 XNOR2_X2 _21978_ (.A(_09809_),
    .B(_09789_),
    .ZN(_12614_));
 XNOR2_X2 _21979_ (.A(_09869_),
    .B(_12614_),
    .ZN(_12615_));
 XNOR2_X1 _21980_ (.A(_09808_),
    .B(_09814_),
    .ZN(_12616_));
 XNOR2_X1 _21981_ (.A(_12615_),
    .B(_12616_),
    .ZN(_12617_));
 MUX2_X2 _21982_ (.A(\text_in_r[85] ),
    .B(_12617_),
    .S(net594),
    .Z(_12618_));
 XOR2_X2 _21983_ (.A(_06270_),
    .B(_12618_),
    .Z(_12619_));
 BUF_X4 _21984_ (.A(_12619_),
    .Z(_12620_));
 BUF_X4 _21985_ (.A(_12620_),
    .Z(_12621_));
 CLKBUF_X3 _21986_ (.A(_12621_),
    .Z(_12622_));
 XNOR2_X2 _21987_ (.A(_09799_),
    .B(_09712_),
    .ZN(_12623_));
 XNOR2_X1 _21988_ (.A(_09788_),
    .B(_12623_),
    .ZN(_12624_));
 XNOR2_X1 _21989_ (.A(_09796_),
    .B(_12624_),
    .ZN(_12625_));
 MUX2_X2 _21990_ (.A(\text_in_r[87] ),
    .B(_12625_),
    .S(_09803_),
    .Z(_12626_));
 XOR2_X2 _21991_ (.A(_06588_),
    .B(_12626_),
    .Z(_12627_));
 XNOR2_X2 _21992_ (.A(_09790_),
    .B(_09798_),
    .ZN(_12628_));
 XNOR2_X2 _21993_ (.A(_09814_),
    .B(_12628_),
    .ZN(_12629_));
 XNOR2_X1 _21994_ (.A(_09785_),
    .B(_09787_),
    .ZN(_12630_));
 XNOR2_X1 _21995_ (.A(_12629_),
    .B(_12630_),
    .ZN(_12631_));
 MUX2_X2 _21996_ (.A(\text_in_r[86] ),
    .B(_12631_),
    .S(_11192_),
    .Z(_12632_));
 XNOR2_X2 _21997_ (.A(_06576_),
    .B(_12632_),
    .ZN(_12633_));
 BUF_X4 _21998_ (.A(_12633_),
    .Z(_12634_));
 NOR3_X1 _21999_ (.A1(_12622_),
    .A2(_12627_),
    .A3(_12634_),
    .ZN(_12635_));
 XNOR2_X2 _22000_ (.A(_06270_),
    .B(_12618_),
    .ZN(_12636_));
 BUF_X4 _22001_ (.A(_12636_),
    .Z(_12637_));
 NAND2_X1 _22002_ (.A1(_12637_),
    .A2(_12633_),
    .ZN(_12638_));
 NOR2_X1 _22003_ (.A1(_12627_),
    .A2(_12638_),
    .ZN(_12639_));
 NOR2_X1 _22004_ (.A1(_12508_),
    .A2(_12543_),
    .ZN(_12640_));
 CLKBUF_X2 split166 (.A(_14874_),
    .Z(net166));
 NAND3_X2 _22006_ (.A1(net203),
    .A2(_12602_),
    .A3(_12603_),
    .ZN(_12642_));
 INV_X8 _22007_ (.A(net500),
    .ZN(_12643_));
 BUF_X4 _22008_ (.A(_12544_),
    .Z(_12644_));
 BUF_X4 _22009_ (.A(_12644_),
    .Z(_12645_));
 NAND2_X1 _22010_ (.A1(_12643_),
    .A2(_12645_),
    .ZN(_12646_));
 OAI22_X1 _22011_ (.A1(_12640_),
    .A2(_12642_),
    .B1(_12646_),
    .B2(_12583_),
    .ZN(_12647_));
 AND2_X2 clone140 (.A1(net546),
    .A2(_12505_),
    .ZN(net140));
 INV_X2 _22013_ (.A(_14964_),
    .ZN(_12649_));
 NAND2_X1 _22014_ (.A1(_12649_),
    .A2(_12607_),
    .ZN(_12650_));
 NOR3_X2 _22015_ (.A1(_12544_),
    .A2(_12586_),
    .A3(_12590_),
    .ZN(_12651_));
 NOR2_X2 _22016_ (.A1(_12598_),
    .A2(_12651_),
    .ZN(_12652_));
 BUF_X8 clone171 (.A(_04387_),
    .Z(net171));
 BUF_X4 _22018_ (.A(_12586_),
    .Z(_12654_));
 BUF_X4 _22019_ (.A(_12590_),
    .Z(_12655_));
 OAI21_X4 _22020_ (.A(_12601_),
    .B1(_12654_),
    .B2(_12655_),
    .ZN(_12656_));
 OAI221_X1 _22021_ (.A(_12650_),
    .B1(_12652_),
    .B2(_14956_),
    .C1(_12656_),
    .C2(_12643_),
    .ZN(_12657_));
 NOR2_X4 _22022_ (.A1(_12561_),
    .A2(_12564_),
    .ZN(_12658_));
 BUF_X4 _22023_ (.A(_12658_),
    .Z(_12659_));
 BUF_X4 _22024_ (.A(_12659_),
    .Z(_12660_));
 BUF_X4 _22025_ (.A(_12660_),
    .Z(_12661_));
 MUX2_X1 _22026_ (.A(_12647_),
    .B(_12657_),
    .S(_12661_),
    .Z(_12662_));
 AOI22_X2 _22027_ (.A1(_12613_),
    .A2(_12635_),
    .B1(_12639_),
    .B2(_12662_),
    .ZN(_12663_));
 XNOR2_X2 _22028_ (.A(_06588_),
    .B(_12626_),
    .ZN(_12664_));
 XOR2_X2 _22029_ (.A(_06576_),
    .B(_12632_),
    .Z(_12665_));
 CLKBUF_X3 _22030_ (.A(_12665_),
    .Z(_12666_));
 BUF_X4 _22031_ (.A(_12660_),
    .Z(_12667_));
 NOR3_X4 _22032_ (.A1(net607),
    .A2(_12586_),
    .A3(_12590_),
    .ZN(_12668_));
 AOI21_X2 _22033_ (.A(net931),
    .B1(_12602_),
    .B2(_12603_),
    .ZN(_12669_));
 AOI21_X2 _22034_ (.A(_12669_),
    .B1(_12592_),
    .B2(net722),
    .ZN(_12670_));
 BUF_X4 rebuffer398 (.A(_04519_),
    .Z(net914));
 AOI221_X1 _22036_ (.A(_12668_),
    .B1(_12670_),
    .B2(_12546_),
    .C1(net202),
    .C2(_12609_),
    .ZN(_12672_));
 NOR2_X2 _22037_ (.A1(_12508_),
    .A2(_12591_),
    .ZN(_12673_));
 NOR2_X1 _22038_ (.A1(_12584_),
    .A2(_12673_),
    .ZN(_12674_));
 BUF_X4 _22039_ (.A(_14961_),
    .Z(_12675_));
 BUF_X8 _22040_ (.A(_12675_),
    .Z(_12676_));
 OAI21_X1 _22041_ (.A(_12661_),
    .B1(_12656_),
    .B2(_12676_),
    .ZN(_12677_));
 OAI221_X1 _22042_ (.A(_12666_),
    .B1(_12667_),
    .B2(_12672_),
    .C1(_12674_),
    .C2(_12677_),
    .ZN(_12678_));
 BUF_X4 _22043_ (.A(_12567_),
    .Z(_12679_));
 NOR2_X1 _22044_ (.A1(_12665_),
    .A2(_12679_),
    .ZN(_12680_));
 BUF_X4 _22045_ (.A(_12644_),
    .Z(_12681_));
 CLKBUF_X3 _22046_ (.A(_12681_),
    .Z(_12682_));
 NOR3_X4 _22047_ (.A1(_12654_),
    .A2(net499),
    .A3(_12655_),
    .ZN(_12683_));
 AOI21_X4 _22048_ (.A(_12649_),
    .B1(_12596_),
    .B2(_12597_),
    .ZN(_12684_));
 NOR3_X1 _22049_ (.A1(_12682_),
    .A2(net911),
    .A3(_12684_),
    .ZN(_12685_));
 BUF_X4 _22050_ (.A(_12601_),
    .Z(_12686_));
 CLKBUF_X3 _22051_ (.A(_12686_),
    .Z(_12687_));
 CLKBUF_X3 _22052_ (.A(_12582_),
    .Z(_12688_));
 BUF_X4 _22053_ (.A(_12688_),
    .Z(_12689_));
 AOI21_X1 _22054_ (.A(_12687_),
    .B1(_12689_),
    .B2(net538),
    .ZN(_12690_));
 NAND2_X4 _22055_ (.A1(_12508_),
    .A2(_12668_),
    .ZN(_12691_));
 AOI21_X1 _22056_ (.A(_12685_),
    .B1(_12690_),
    .B2(_12691_),
    .ZN(_12692_));
 NOR2_X2 _22057_ (.A1(_12665_),
    .A2(_12660_),
    .ZN(_12693_));
 NOR2_X2 _22058_ (.A1(_12548_),
    .A2(_12545_),
    .ZN(_12694_));
 BUF_X4 _22059_ (.A(_12606_),
    .Z(_12695_));
 AOI21_X1 _22060_ (.A(_12694_),
    .B1(_14954_),
    .B2(_12695_),
    .ZN(_12696_));
 XNOR2_X1 _22061_ (.A(_12689_),
    .B(_12696_),
    .ZN(_12697_));
 AOI22_X1 _22062_ (.A1(_12680_),
    .A2(_12692_),
    .B1(_12693_),
    .B2(_12697_),
    .ZN(_12698_));
 NAND4_X1 _22063_ (.A1(_12622_),
    .A2(_12664_),
    .A3(_12678_),
    .A4(_12698_),
    .ZN(_12699_));
 NOR2_X2 _22064_ (.A1(_12636_),
    .A2(_12665_),
    .ZN(_12700_));
 CLKBUF_X3 _22065_ (.A(_12581_),
    .Z(_12701_));
 CLKBUF_X3 _22066_ (.A(_12701_),
    .Z(_12702_));
 OAI21_X4 _22067_ (.A(_12548_),
    .B1(_12586_),
    .B2(_12590_),
    .ZN(_12703_));
 OAI221_X1 _22068_ (.A(_12687_),
    .B1(_12702_),
    .B2(_12605_),
    .C1(_12703_),
    .C2(net200),
    .ZN(_12704_));
 BUF_X8 _22069_ (.A(_14966_),
    .Z(_12705_));
 NAND2_X1 _22070_ (.A1(_12705_),
    .A2(_12599_),
    .ZN(_12706_));
 AND3_X1 _22071_ (.A1(_12667_),
    .A2(_12704_),
    .A3(_12706_),
    .ZN(_12707_));
 NAND3_X4 _22072_ (.A1(_12545_),
    .A2(_12602_),
    .A3(_12603_),
    .ZN(_12708_));
 NOR2_X1 _22073_ (.A1(_14964_),
    .A2(_12708_),
    .ZN(_12709_));
 INV_X1 _22074_ (.A(_12605_),
    .ZN(_12710_));
 NOR3_X4 _22075_ (.A1(_12527_),
    .A2(_12654_),
    .A3(_12655_),
    .ZN(_12711_));
 AOI221_X2 _22076_ (.A(_12546_),
    .B1(_12582_),
    .B2(_12710_),
    .C1(_12711_),
    .C2(net723),
    .ZN(_12712_));
 NOR3_X1 _22077_ (.A1(_12667_),
    .A2(_12709_),
    .A3(_12712_),
    .ZN(_12713_));
 OAI21_X1 _22078_ (.A(_12700_),
    .B1(_12707_),
    .B2(_12713_),
    .ZN(_12714_));
 CLKBUF_X3 _22079_ (.A(_12637_),
    .Z(_12715_));
 BUF_X4 _22080_ (.A(_12715_),
    .Z(_12716_));
 NOR2_X1 _22081_ (.A1(_12716_),
    .A2(_12634_),
    .ZN(_12717_));
 NOR3_X4 _22082_ (.A1(_12605_),
    .A2(_12654_),
    .A3(_12655_),
    .ZN(_12718_));
 AOI21_X4 _22083_ (.A(_12676_),
    .B1(_12602_),
    .B2(_12603_),
    .ZN(_12719_));
 NOR2_X1 _22084_ (.A1(_12718_),
    .A2(_12719_),
    .ZN(_12720_));
 NOR2_X1 _22085_ (.A1(_14979_),
    .A2(_12720_),
    .ZN(_12721_));
 INV_X2 _22086_ (.A(_14956_),
    .ZN(_12722_));
 OAI21_X1 _22087_ (.A(_12568_),
    .B1(_12708_),
    .B2(_12722_),
    .ZN(_12723_));
 AOI21_X4 _22088_ (.A(net608),
    .B1(_12596_),
    .B2(_12597_),
    .ZN(_12724_));
 BUF_X4 _22089_ (.A(_12591_),
    .Z(_12725_));
 CLKBUF_X3 _22090_ (.A(_12725_),
    .Z(_12726_));
 AOI21_X1 _22091_ (.A(_12724_),
    .B1(_12726_),
    .B2(_14955_),
    .ZN(_12727_));
 AOI21_X2 _22092_ (.A(_12683_),
    .B1(_12702_),
    .B2(_12649_),
    .ZN(_12728_));
 MUX2_X1 _22093_ (.A(_12727_),
    .B(_12728_),
    .S(_12682_),
    .Z(_12729_));
 OAI221_X2 _22094_ (.A(_12717_),
    .B1(_12721_),
    .B2(_12723_),
    .C1(_12612_),
    .C2(_12729_),
    .ZN(_12730_));
 NAND3_X2 _22095_ (.A1(_12627_),
    .A2(_12730_),
    .A3(_12714_),
    .ZN(_12731_));
 AOI21_X4 _22096_ (.A(net501),
    .B1(_12596_),
    .B2(_12597_),
    .ZN(_12732_));
 NOR3_X2 _22097_ (.A1(_12705_),
    .A2(_12654_),
    .A3(_12655_),
    .ZN(_12733_));
 OAI21_X1 _22098_ (.A(_12687_),
    .B1(_12732_),
    .B2(_12733_),
    .ZN(_12734_));
 INV_X2 _22099_ (.A(_12675_),
    .ZN(_12735_));
 NAND2_X1 _22100_ (.A1(_12735_),
    .A2(_12607_),
    .ZN(_12736_));
 NAND4_X1 _22101_ (.A1(_12666_),
    .A2(_12568_),
    .A3(_12734_),
    .A4(_12736_),
    .ZN(_12737_));
 NAND2_X1 _22102_ (.A1(_12735_),
    .A2(_12726_),
    .ZN(_12738_));
 NAND4_X1 _22103_ (.A1(_12665_),
    .A2(_12661_),
    .A3(_12600_),
    .A4(_12738_),
    .ZN(_12739_));
 AOI21_X4 _22104_ (.A(_12548_),
    .B1(_12505_),
    .B2(net546),
    .ZN(_12740_));
 NOR2_X2 _22105_ (.A1(_12592_),
    .A2(_12740_),
    .ZN(_12741_));
 NOR2_X1 _22106_ (.A1(_14979_),
    .A2(_12741_),
    .ZN(_12742_));
 OAI21_X1 _22107_ (.A(_12737_),
    .B1(_12739_),
    .B2(_12742_),
    .ZN(_12743_));
 NAND2_X1 _22108_ (.A1(net502),
    .A2(_12545_),
    .ZN(_12744_));
 NAND2_X1 _22109_ (.A1(_12592_),
    .A2(_12744_),
    .ZN(_12745_));
 OAI21_X1 _22110_ (.A(_12745_),
    .B1(_12725_),
    .B2(_14977_),
    .ZN(_12746_));
 NOR2_X2 _22111_ (.A1(_12527_),
    .A2(_12544_),
    .ZN(_12747_));
 AOI22_X4 _22112_ (.A1(_12735_),
    .A2(_12545_),
    .B1(_12747_),
    .B2(net722),
    .ZN(_12748_));
 AOI21_X4 _22113_ (.A(_12566_),
    .B1(_12592_),
    .B2(_12748_),
    .ZN(_12749_));
 NAND3_X2 _22114_ (.A1(_12605_),
    .A2(_12602_),
    .A3(_12603_),
    .ZN(_12750_));
 OAI21_X4 _22115_ (.A(_12527_),
    .B1(_12586_),
    .B2(_12590_),
    .ZN(_12751_));
 AOI21_X1 _22116_ (.A(_12551_),
    .B1(_12750_),
    .B2(_12751_),
    .ZN(_12752_));
 AOI21_X1 _22117_ (.A(_12752_),
    .B1(_12609_),
    .B2(_12722_),
    .ZN(_12753_));
 AOI221_X2 _22118_ (.A(_12665_),
    .B1(_12679_),
    .B2(_12746_),
    .C1(_12749_),
    .C2(_12753_),
    .ZN(_12754_));
 NOR3_X1 _22119_ (.A1(_12622_),
    .A2(_12743_),
    .A3(_12754_),
    .ZN(_12755_));
 OAI211_X2 _22120_ (.A(_12663_),
    .B(_12699_),
    .C1(_12755_),
    .C2(_12731_),
    .ZN(_00072_));
 NAND2_X1 _22121_ (.A1(_12664_),
    .A2(_12665_),
    .ZN(_12756_));
 BUF_X4 _22122_ (.A(_12620_),
    .Z(_12757_));
 NAND2_X1 _22123_ (.A1(_12701_),
    .A2(_12740_),
    .ZN(_12758_));
 NOR2_X1 _22124_ (.A1(_12551_),
    .A2(_12718_),
    .ZN(_12759_));
 NOR3_X4 _22125_ (.A1(_12590_),
    .A2(_12586_),
    .A3(_14970_),
    .ZN(_12760_));
 NOR2_X1 _22126_ (.A1(_12681_),
    .A2(_12760_),
    .ZN(_12761_));
 OAI21_X4 _22127_ (.A(net501),
    .B1(_12654_),
    .B2(_12655_),
    .ZN(_12762_));
 AOI221_X2 _22128_ (.A(_12757_),
    .B1(_12758_),
    .B2(_12759_),
    .C1(_12761_),
    .C2(_12762_),
    .ZN(_12763_));
 NOR3_X2 _22129_ (.A1(_12686_),
    .A2(_12711_),
    .A3(net673),
    .ZN(_12764_));
 OAI21_X2 _22130_ (.A(_12722_),
    .B1(_12654_),
    .B2(_12655_),
    .ZN(_12765_));
 AOI21_X1 _22131_ (.A(_12547_),
    .B1(_12750_),
    .B2(_12765_),
    .ZN(_12766_));
 NOR3_X1 _22132_ (.A1(_12716_),
    .A2(_12764_),
    .A3(_12766_),
    .ZN(_12767_));
 OAI21_X1 _22133_ (.A(_12612_),
    .B1(_12763_),
    .B2(_12767_),
    .ZN(_12768_));
 OAI21_X2 _22134_ (.A(_12643_),
    .B1(_12654_),
    .B2(_12655_),
    .ZN(_12769_));
 AOI21_X1 _22135_ (.A(_12682_),
    .B1(_12769_),
    .B2(_12691_),
    .ZN(_12770_));
 OAI21_X1 _22136_ (.A(_12715_),
    .B1(_12708_),
    .B2(_14963_),
    .ZN(_12771_));
 NAND3_X4 _22137_ (.A1(_12548_),
    .A2(_12602_),
    .A3(_12603_),
    .ZN(_12772_));
 OAI21_X1 _22138_ (.A(_12676_),
    .B1(_12654_),
    .B2(_12655_),
    .ZN(_12773_));
 AOI21_X2 _22139_ (.A(_12645_),
    .B1(_12772_),
    .B2(_12773_),
    .ZN(_12774_));
 BUF_X4 _22140_ (.A(_12508_),
    .Z(_12775_));
 MUX2_X1 _22141_ (.A(_12722_),
    .B(_12775_),
    .S(_12688_),
    .Z(_12776_));
 AOI21_X1 _22142_ (.A(_12774_),
    .B1(_12776_),
    .B2(_14979_),
    .ZN(_12777_));
 OAI221_X1 _22143_ (.A(_12667_),
    .B1(_12770_),
    .B2(_12771_),
    .C1(_12777_),
    .C2(_12716_),
    .ZN(_12778_));
 AOI21_X1 _22144_ (.A(_12756_),
    .B1(_12768_),
    .B2(_12778_),
    .ZN(_12779_));
 NOR2_X2 _22145_ (.A1(_12664_),
    .A2(_12634_),
    .ZN(_12780_));
 BUF_X4 _22146_ (.A(_12651_),
    .Z(_12781_));
 OAI21_X1 _22147_ (.A(_14954_),
    .B1(_12599_),
    .B2(_12781_),
    .ZN(_12782_));
 AOI22_X1 _22148_ (.A1(net202),
    .A2(_12607_),
    .B1(_12724_),
    .B2(net200),
    .ZN(_12783_));
 NAND3_X1 _22149_ (.A1(_12716_),
    .A2(_12782_),
    .A3(_12783_),
    .ZN(_12784_));
 OAI21_X1 _22150_ (.A(_12547_),
    .B1(_12726_),
    .B2(_12740_),
    .ZN(_12785_));
 NAND3_X4 _22151_ (.A1(_12675_),
    .A2(_12596_),
    .A3(_12597_),
    .ZN(_12786_));
 NAND3_X1 _22152_ (.A1(_12687_),
    .A2(_12769_),
    .A3(_12786_),
    .ZN(_12787_));
 NAND3_X1 _22153_ (.A1(_12621_),
    .A2(_12785_),
    .A3(_12787_),
    .ZN(_12788_));
 NAND4_X1 _22154_ (.A1(_12667_),
    .A2(_12780_),
    .A3(_12784_),
    .A4(_12788_),
    .ZN(_12789_));
 NAND2_X1 _22155_ (.A1(_12612_),
    .A2(_12780_),
    .ZN(_12790_));
 INV_X4 _22156_ (.A(net931),
    .ZN(_12791_));
 AOI21_X4 _22157_ (.A(_12791_),
    .B1(_12602_),
    .B2(_12603_),
    .ZN(_12792_));
 NOR2_X1 _22158_ (.A1(_14972_),
    .A2(_12792_),
    .ZN(_12793_));
 NOR2_X1 _22159_ (.A1(_14960_),
    .A2(_12656_),
    .ZN(_12794_));
 NAND2_X1 _22160_ (.A1(_12621_),
    .A2(_12691_),
    .ZN(_12795_));
 NOR3_X4 _22161_ (.A1(_12722_),
    .A2(_12586_),
    .A3(_12590_),
    .ZN(_12796_));
 AOI21_X2 _22162_ (.A(_12643_),
    .B1(_12596_),
    .B2(_12597_),
    .ZN(_12797_));
 NOR2_X2 _22163_ (.A1(_12797_),
    .A2(_12796_),
    .ZN(_12798_));
 NOR2_X1 _22164_ (.A1(_12547_),
    .A2(_12798_),
    .ZN(_12799_));
 NOR2_X1 _22165_ (.A1(_12735_),
    .A2(_12725_),
    .ZN(_12800_));
 NOR3_X1 _22166_ (.A1(_12552_),
    .A2(_12800_),
    .A3(_12668_),
    .ZN(_12801_));
 OAI33_X1 _22167_ (.A1(_12793_),
    .A2(_12794_),
    .A3(_12795_),
    .B1(_12799_),
    .B2(_12801_),
    .B3(_12621_),
    .ZN(_12802_));
 OAI21_X1 _22168_ (.A(_12789_),
    .B1(_12802_),
    .B2(_12790_),
    .ZN(_12803_));
 OAI21_X1 _22169_ (.A(_12744_),
    .B1(_12644_),
    .B2(_12791_),
    .ZN(_12804_));
 NAND2_X1 _22170_ (.A1(_12701_),
    .A2(_12804_),
    .ZN(_12805_));
 OAI21_X1 _22171_ (.A(_12736_),
    .B1(_12652_),
    .B2(_12695_),
    .ZN(_12806_));
 AOI221_X2 _22172_ (.A(_12757_),
    .B1(_12805_),
    .B2(_12749_),
    .C1(_12806_),
    .C2(_12679_),
    .ZN(_12807_));
 NAND2_X2 _22173_ (.A1(_12566_),
    .A2(_12591_),
    .ZN(_12808_));
 MUX2_X1 _22174_ (.A(_12675_),
    .B(_12548_),
    .S(_12545_),
    .Z(_12809_));
 NOR2_X1 _22175_ (.A1(_12643_),
    .A2(_12659_),
    .ZN(_12810_));
 OAI221_X2 _22176_ (.A(_12620_),
    .B1(_12808_),
    .B2(_12809_),
    .C1(_12810_),
    .C2(_12656_),
    .ZN(_12811_));
 NAND3_X1 _22177_ (.A1(_12644_),
    .A2(_12566_),
    .A3(_12582_),
    .ZN(_12812_));
 NAND3_X1 _22178_ (.A1(net139),
    .A2(_12659_),
    .A3(_12592_),
    .ZN(_12813_));
 NAND2_X1 _22179_ (.A1(_12812_),
    .A2(_12813_),
    .ZN(_12814_));
 OAI21_X1 _22180_ (.A(_12600_),
    .B1(_12567_),
    .B2(_12645_),
    .ZN(_12815_));
 AOI221_X2 _22181_ (.A(_12811_),
    .B1(_12814_),
    .B2(_12549_),
    .C1(_12815_),
    .C2(_14960_),
    .ZN(_12816_));
 NAND2_X2 _22182_ (.A1(_12627_),
    .A2(_12634_),
    .ZN(_12817_));
 NOR3_X2 _22183_ (.A1(_12807_),
    .A2(_12816_),
    .A3(_12817_),
    .ZN(_12818_));
 NAND2_X1 _22184_ (.A1(_12664_),
    .A2(_12634_),
    .ZN(_12819_));
 NAND2_X1 _22185_ (.A1(_12508_),
    .A2(_12582_),
    .ZN(_12820_));
 XNOR2_X2 _22186_ (.A(_12527_),
    .B(_12546_),
    .ZN(_12821_));
 AOI21_X1 _22187_ (.A(_12747_),
    .B1(_12681_),
    .B2(_14956_),
    .ZN(_12822_));
 OAI221_X1 _22188_ (.A(_12757_),
    .B1(_12820_),
    .B2(_12821_),
    .C1(_12822_),
    .C2(_12702_),
    .ZN(_12823_));
 XNOR2_X1 _22189_ (.A(_12695_),
    .B(_12725_),
    .ZN(_12824_));
 AOI21_X1 _22190_ (.A(_12774_),
    .B1(_12824_),
    .B2(_12682_),
    .ZN(_12825_));
 OAI221_X1 _22191_ (.A(_12823_),
    .B1(_12564_),
    .B2(_12561_),
    .C1(_12825_),
    .C2(_12621_),
    .ZN(_12826_));
 MUX2_X1 _22192_ (.A(_14964_),
    .B(_12740_),
    .S(_12550_),
    .Z(_12827_));
 NAND2_X1 _22193_ (.A1(_12636_),
    .A2(_12581_),
    .ZN(_12828_));
 OAI221_X2 _22194_ (.A(_12661_),
    .B1(_12689_),
    .B2(_12827_),
    .C1(_12828_),
    .C2(_14980_),
    .ZN(_12829_));
 AOI21_X2 _22195_ (.A(_12819_),
    .B1(_12826_),
    .B2(_12829_),
    .ZN(_12830_));
 NOR4_X2 _22196_ (.A1(_12779_),
    .A2(_12803_),
    .A3(_12818_),
    .A4(_12830_),
    .ZN(_00073_));
 NAND2_X1 _22197_ (.A1(_12642_),
    .A2(_12751_),
    .ZN(_12831_));
 MUX2_X1 _22198_ (.A(_12605_),
    .B(_12606_),
    .S(_12591_),
    .Z(_12832_));
 MUX2_X1 _22199_ (.A(_12831_),
    .B(_12832_),
    .S(_12546_),
    .Z(_12833_));
 NOR2_X2 _22200_ (.A1(_12637_),
    .A2(_12659_),
    .ZN(_12834_));
 AND2_X1 _22201_ (.A1(_12833_),
    .A2(_12834_),
    .ZN(_12835_));
 INV_X1 _22202_ (.A(_12819_),
    .ZN(_12836_));
 NAND2_X2 _22203_ (.A1(_12620_),
    .A2(_12658_),
    .ZN(_12837_));
 AOI21_X2 _22204_ (.A(_12527_),
    .B1(_12602_),
    .B2(_12603_),
    .ZN(_12838_));
 OR4_X1 _22205_ (.A1(net139),
    .A2(_12601_),
    .A3(_12838_),
    .A4(_12668_),
    .ZN(_12839_));
 OAI21_X1 _22206_ (.A(_12839_),
    .B1(_12656_),
    .B2(net138),
    .ZN(_12840_));
 OAI21_X1 _22207_ (.A(_12836_),
    .B1(_12837_),
    .B2(_12840_),
    .ZN(_12841_));
 NOR2_X4 _22208_ (.A1(_12619_),
    .A2(_12566_),
    .ZN(_12842_));
 NOR2_X1 _22209_ (.A1(_12695_),
    .A2(_12546_),
    .ZN(_12843_));
 OAI221_X1 _22210_ (.A(_12842_),
    .B1(_12843_),
    .B2(_12745_),
    .C1(_12593_),
    .C2(_12748_),
    .ZN(_12844_));
 NAND2_X1 _22211_ (.A1(_12637_),
    .A2(_12679_),
    .ZN(_12845_));
 NAND3_X2 _22212_ (.A1(net931),
    .A2(_12596_),
    .A3(_12597_),
    .ZN(_12846_));
 NAND2_X1 _22213_ (.A1(_12751_),
    .A2(_12846_),
    .ZN(_12847_));
 AOI221_X1 _22214_ (.A(_12673_),
    .B1(_12847_),
    .B2(_12644_),
    .C1(_12781_),
    .C2(_12676_),
    .ZN(_12848_));
 OAI21_X1 _22215_ (.A(_12844_),
    .B1(_12845_),
    .B2(_12848_),
    .ZN(_12849_));
 NOR2_X4 _22216_ (.A1(_12620_),
    .A2(_12658_),
    .ZN(_12850_));
 OR2_X4 _22217_ (.A1(_12550_),
    .A2(_12760_),
    .ZN(_12851_));
 OR2_X1 _22218_ (.A1(_12838_),
    .A2(_12733_),
    .ZN(_12852_));
 OAI22_X1 _22219_ (.A1(_12719_),
    .A2(_12851_),
    .B1(_12852_),
    .B2(_12645_),
    .ZN(_12853_));
 AND2_X1 _22220_ (.A1(_12850_),
    .A2(_12853_),
    .ZN(_12854_));
 NOR2_X2 _22221_ (.A1(_12627_),
    .A2(_12634_),
    .ZN(_12855_));
 INV_X16 _22222_ (.A(_12705_),
    .ZN(_12856_));
 OAI21_X1 _22223_ (.A(_12551_),
    .B1(_12582_),
    .B2(_12856_),
    .ZN(_12857_));
 NOR2_X2 _22224_ (.A1(_12606_),
    .A2(_12591_),
    .ZN(_12858_));
 OAI221_X1 _22225_ (.A(_12842_),
    .B1(_12857_),
    .B2(_12858_),
    .C1(_12686_),
    .C2(_12676_),
    .ZN(_12859_));
 BUF_X4 _22226_ (.A(_12658_),
    .Z(_12860_));
 OAI21_X1 _22227_ (.A(_12551_),
    .B1(_12711_),
    .B2(_12732_),
    .ZN(_12861_));
 OAI21_X1 _22228_ (.A(_12644_),
    .B1(_12733_),
    .B2(_12797_),
    .ZN(_12862_));
 NAND4_X1 _22229_ (.A1(_12862_),
    .A2(_12860_),
    .A3(_12861_),
    .A4(_12620_),
    .ZN(_12863_));
 NAND3_X1 _22230_ (.A1(_12855_),
    .A2(_12859_),
    .A3(_12863_),
    .ZN(_12864_));
 OAI21_X1 _22231_ (.A(_12772_),
    .B1(_12592_),
    .B2(_12705_),
    .ZN(_12865_));
 OAI22_X1 _22232_ (.A1(_12645_),
    .A2(_12865_),
    .B1(_12851_),
    .B2(_12858_),
    .ZN(_12866_));
 AND2_X1 _22233_ (.A1(_12834_),
    .A2(_12866_),
    .ZN(_12867_));
 OAI33_X1 _22234_ (.A1(_12835_),
    .A2(_12841_),
    .A3(_12849_),
    .B1(_12864_),
    .B2(_12854_),
    .B3(_12867_),
    .ZN(_12868_));
 NAND2_X1 _22235_ (.A1(_14977_),
    .A2(_12592_),
    .ZN(_12869_));
 NAND2_X1 _22236_ (.A1(_12548_),
    .A2(_12550_),
    .ZN(_12870_));
 OAI221_X2 _22237_ (.A(_12582_),
    .B1(_12870_),
    .B2(net139),
    .C1(_12601_),
    .C2(net499),
    .ZN(_12871_));
 AOI21_X1 _22238_ (.A(_12837_),
    .B1(_12869_),
    .B2(_12871_),
    .ZN(_12872_));
 AOI21_X1 _22239_ (.A(_12684_),
    .B1(_12591_),
    .B2(_12506_),
    .ZN(_12873_));
 NOR2_X2 _22240_ (.A1(_12732_),
    .A2(_12796_),
    .ZN(_12874_));
 MUX2_X1 _22241_ (.A(_12873_),
    .B(_12874_),
    .S(_12545_),
    .Z(_12875_));
 AND2_X1 _22242_ (.A1(_14980_),
    .A2(_12591_),
    .ZN(_12876_));
 MUX2_X1 _22243_ (.A(_12548_),
    .B(_12550_),
    .S(_12508_),
    .Z(_12877_));
 AOI21_X1 _22244_ (.A(_12876_),
    .B1(_12877_),
    .B2(_12581_),
    .ZN(_12878_));
 MUX2_X1 _22245_ (.A(_12875_),
    .B(_12878_),
    .S(_12658_),
    .Z(_12879_));
 NOR3_X1 _22246_ (.A1(net140),
    .A2(_12545_),
    .A3(_12724_),
    .ZN(_12880_));
 NAND2_X2 _22247_ (.A1(_12527_),
    .A2(_12550_),
    .ZN(_12881_));
 NOR2_X2 _22248_ (.A1(_12506_),
    .A2(_12581_),
    .ZN(_12882_));
 OR2_X1 _22249_ (.A1(_12882_),
    .A2(_12640_),
    .ZN(_12883_));
 AOI221_X2 _22250_ (.A(_12880_),
    .B1(_12881_),
    .B2(_12673_),
    .C1(net202),
    .C2(_12883_),
    .ZN(_12884_));
 AOI221_X2 _22251_ (.A(_12872_),
    .B1(_12879_),
    .B2(_12637_),
    .C1(_12834_),
    .C2(_12884_),
    .ZN(_12885_));
 AOI21_X1 _22252_ (.A(_12820_),
    .B1(_12547_),
    .B2(_14963_),
    .ZN(_12886_));
 OAI21_X1 _22253_ (.A(_12715_),
    .B1(_12702_),
    .B2(_14984_),
    .ZN(_12887_));
 NOR2_X1 _22254_ (.A1(_12688_),
    .A2(_12740_),
    .ZN(_12888_));
 NOR2_X2 _22255_ (.A1(_14958_),
    .A2(_12675_),
    .ZN(_12889_));
 OAI21_X1 _22256_ (.A(_12552_),
    .B1(_12593_),
    .B2(_12889_),
    .ZN(_12890_));
 NAND3_X2 _22257_ (.A1(_12649_),
    .A2(_12602_),
    .A3(_12603_),
    .ZN(_12891_));
 NAND2_X1 _22258_ (.A1(_12681_),
    .A2(_12891_),
    .ZN(_12892_));
 OAI22_X1 _22259_ (.A1(_12888_),
    .A2(_12890_),
    .B1(_12892_),
    .B2(_12741_),
    .ZN(_12893_));
 OAI221_X2 _22260_ (.A(_12568_),
    .B1(_12886_),
    .B2(_12887_),
    .C1(_12893_),
    .C2(_12716_),
    .ZN(_12894_));
 AOI21_X1 _22261_ (.A(_12527_),
    .B1(_12505_),
    .B2(net548),
    .ZN(_12895_));
 NAND3_X1 _22262_ (.A1(_12681_),
    .A2(_12593_),
    .A3(_12895_),
    .ZN(_12896_));
 NAND2_X1 _22263_ (.A1(_14975_),
    .A2(_12688_),
    .ZN(_12897_));
 AOI21_X1 _22264_ (.A(_12757_),
    .B1(_12896_),
    .B2(_12897_),
    .ZN(_12898_));
 AOI22_X1 _22265_ (.A1(_12676_),
    .A2(_12599_),
    .B1(_12874_),
    .B2(_12687_),
    .ZN(_12899_));
 AOI21_X1 _22266_ (.A(_12898_),
    .B1(_12899_),
    .B2(_12621_),
    .ZN(_12900_));
 OAI21_X2 _22267_ (.A(_12894_),
    .B1(_12900_),
    .B2(_12612_),
    .ZN(_12901_));
 INV_X1 _22268_ (.A(_12817_),
    .ZN(_12902_));
 AOI221_X1 _22269_ (.A(_12868_),
    .B1(_12780_),
    .B2(_12885_),
    .C1(_12901_),
    .C2(_12902_),
    .ZN(_00074_));
 INV_X1 _22270_ (.A(_12780_),
    .ZN(_12903_));
 NOR2_X4 _22271_ (.A1(net140),
    .A2(_12703_),
    .ZN(_12904_));
 AOI21_X1 _22272_ (.A(_12687_),
    .B1(_12751_),
    .B2(_12891_),
    .ZN(_12905_));
 NOR2_X1 _22273_ (.A1(net499),
    .A2(_12604_),
    .ZN(_12906_));
 NOR3_X1 _22274_ (.A1(_12904_),
    .A2(_12905_),
    .A3(_12906_),
    .ZN(_12907_));
 AOI21_X1 _22275_ (.A(_12903_),
    .B1(_12834_),
    .B2(_12907_),
    .ZN(_12908_));
 AOI221_X2 _22276_ (.A(_12757_),
    .B1(_12567_),
    .B2(_12906_),
    .C1(_12609_),
    .C2(_12775_),
    .ZN(_12909_));
 AOI21_X1 _22277_ (.A(_12609_),
    .B1(_14954_),
    .B2(net200),
    .ZN(_12910_));
 OAI21_X1 _22278_ (.A(_12909_),
    .B1(_12910_),
    .B2(_12612_),
    .ZN(_12911_));
 NAND2_X1 _22279_ (.A1(net138),
    .A2(_12701_),
    .ZN(_12912_));
 AOI21_X1 _22280_ (.A(_12860_),
    .B1(_12725_),
    .B2(_12705_),
    .ZN(_12913_));
 AOI221_X2 _22281_ (.A(_12552_),
    .B1(_12912_),
    .B2(_12913_),
    .C1(_12660_),
    .C2(_14954_),
    .ZN(_12914_));
 NAND2_X1 _22282_ (.A1(_12527_),
    .A2(_12781_),
    .ZN(_12915_));
 AOI21_X1 _22283_ (.A(_12695_),
    .B1(_12600_),
    .B2(_12915_),
    .ZN(_12916_));
 AOI221_X2 _22284_ (.A(_12916_),
    .B1(_12609_),
    .B2(net666),
    .C1(_12643_),
    .C2(_12607_),
    .ZN(_12917_));
 OAI221_X1 _22285_ (.A(_12908_),
    .B1(_12911_),
    .B2(_12914_),
    .C1(_12917_),
    .C2(_12837_),
    .ZN(_12918_));
 NAND3_X1 _22286_ (.A1(_12682_),
    .A2(_12769_),
    .A3(_12891_),
    .ZN(_12919_));
 OAI21_X1 _22287_ (.A(_12919_),
    .B1(_12832_),
    .B2(_14979_),
    .ZN(_12920_));
 OAI21_X2 _22288_ (.A(_12681_),
    .B1(_12792_),
    .B2(_12668_),
    .ZN(_12921_));
 NAND2_X1 _22289_ (.A1(_12715_),
    .A2(_12660_),
    .ZN(_12922_));
 NAND2_X1 _22290_ (.A1(_12702_),
    .A2(_12889_),
    .ZN(_12923_));
 NOR2_X1 _22291_ (.A1(_12547_),
    .A2(net911),
    .ZN(_12924_));
 AOI21_X1 _22292_ (.A(_12922_),
    .B1(_12923_),
    .B2(_12924_),
    .ZN(_12925_));
 AOI22_X1 _22293_ (.A1(_12850_),
    .A2(_12920_),
    .B1(_12921_),
    .B2(_12925_),
    .ZN(_12926_));
 NAND2_X1 _22294_ (.A1(_14972_),
    .A2(_12568_),
    .ZN(_12927_));
 AOI21_X1 _22295_ (.A(_12683_),
    .B1(_12689_),
    .B2(_12605_),
    .ZN(_12928_));
 AOI22_X1 _22296_ (.A1(_14963_),
    .A2(_12781_),
    .B1(_12652_),
    .B2(_12705_),
    .ZN(_12929_));
 OAI221_X1 _22297_ (.A(_12622_),
    .B1(_12927_),
    .B2(_12928_),
    .C1(_12929_),
    .C2(_12568_),
    .ZN(_12930_));
 AOI21_X1 _22298_ (.A(_12666_),
    .B1(_12926_),
    .B2(_12930_),
    .ZN(_12931_));
 OR2_X1 _22299_ (.A1(_12701_),
    .A2(_12827_),
    .ZN(_12932_));
 INV_X1 _22300_ (.A(_12889_),
    .ZN(_12933_));
 MUX2_X1 _22301_ (.A(_12705_),
    .B(_12933_),
    .S(_12550_),
    .Z(_12934_));
 AOI21_X1 _22302_ (.A(_12620_),
    .B1(_12701_),
    .B2(_12934_),
    .ZN(_12935_));
 OAI21_X1 _22303_ (.A(_14963_),
    .B1(_12681_),
    .B2(_12583_),
    .ZN(_12936_));
 AOI221_X2 _22304_ (.A(_12637_),
    .B1(_12607_),
    .B2(net722),
    .C1(_12608_),
    .C2(_12722_),
    .ZN(_12937_));
 AOI221_X2 _22305_ (.A(_12679_),
    .B1(_12932_),
    .B2(_12935_),
    .C1(_12936_),
    .C2(_12937_),
    .ZN(_12938_));
 NOR2_X2 _22306_ (.A1(_12645_),
    .A2(_12860_),
    .ZN(_12939_));
 OAI21_X1 _22307_ (.A(_12642_),
    .B1(_12593_),
    .B2(_12856_),
    .ZN(_12940_));
 NAND2_X1 _22308_ (.A1(_12637_),
    .A2(_12593_),
    .ZN(_12941_));
 OAI221_X1 _22309_ (.A(_12939_),
    .B1(_12940_),
    .B2(_12715_),
    .C1(_12941_),
    .C2(_14963_),
    .ZN(_12942_));
 NOR2_X1 _22310_ (.A1(_12552_),
    .A2(_12660_),
    .ZN(_12943_));
 OAI221_X2 _22311_ (.A(_12943_),
    .B1(_12751_),
    .B2(_12715_),
    .C1(net138),
    .C2(_12689_),
    .ZN(_12944_));
 NAND3_X1 _22312_ (.A1(_12666_),
    .A2(_12942_),
    .A3(_12944_),
    .ZN(_12945_));
 OAI21_X1 _22313_ (.A(_12664_),
    .B1(_12938_),
    .B2(_12945_),
    .ZN(_12946_));
 XNOR2_X1 _22314_ (.A(_12547_),
    .B(_12660_),
    .ZN(_12947_));
 NAND2_X1 _22315_ (.A1(_12644_),
    .A2(_12659_),
    .ZN(_12948_));
 OAI221_X1 _22316_ (.A(_12689_),
    .B1(_12947_),
    .B2(net202),
    .C1(_12948_),
    .C2(_14960_),
    .ZN(_12949_));
 NOR4_X2 _22317_ (.A1(net723),
    .A2(_12566_),
    .A3(_12582_),
    .A4(_12694_),
    .ZN(_12950_));
 AOI21_X1 _22318_ (.A(_12551_),
    .B1(_12860_),
    .B2(_12549_),
    .ZN(_12951_));
 AOI221_X2 _22319_ (.A(_12950_),
    .B1(_12951_),
    .B2(_12882_),
    .C1(_14963_),
    .C2(_12939_),
    .ZN(_12952_));
 NAND3_X1 _22320_ (.A1(_12716_),
    .A2(_12949_),
    .A3(_12952_),
    .ZN(_12953_));
 NAND2_X1 _22321_ (.A1(_12765_),
    .A2(_12891_),
    .ZN(_12954_));
 OR2_X1 _22322_ (.A1(net673),
    .A2(_12668_),
    .ZN(_12955_));
 MUX2_X1 _22323_ (.A(_12954_),
    .B(_12955_),
    .S(_12681_),
    .Z(_12956_));
 AOI21_X1 _22324_ (.A(_12669_),
    .B1(_12725_),
    .B2(net499),
    .ZN(_12957_));
 AOI21_X1 _22325_ (.A(_12719_),
    .B1(_12725_),
    .B2(_12695_),
    .ZN(_12958_));
 MUX2_X1 _22326_ (.A(_12957_),
    .B(_12958_),
    .S(_12681_),
    .Z(_12959_));
 MUX2_X1 _22327_ (.A(_12956_),
    .B(_12959_),
    .S(_12661_),
    .Z(_12960_));
 OAI21_X2 _22328_ (.A(_12953_),
    .B1(_12960_),
    .B2(_12716_),
    .ZN(_12961_));
 OAI221_X1 _22329_ (.A(_12918_),
    .B1(_12931_),
    .B2(_12946_),
    .C1(_12961_),
    .C2(_12817_),
    .ZN(_00075_));
 OR2_X4 _22330_ (.A1(_12760_),
    .A2(_12644_),
    .ZN(_12962_));
 NOR3_X4 _22331_ (.A1(_12962_),
    .A2(_12904_),
    .A3(_12567_),
    .ZN(_12963_));
 AND2_X4 _22332_ (.A1(_12786_),
    .A2(_12544_),
    .ZN(_12964_));
 AOI221_X2 _22333_ (.A(_12658_),
    .B1(_12762_),
    .B2(_12964_),
    .C1(_12601_),
    .C2(_12856_),
    .ZN(_12965_));
 AOI21_X4 _22334_ (.A(_12856_),
    .B1(_12596_),
    .B2(_12597_),
    .ZN(_12966_));
 AOI21_X4 _22335_ (.A(_12966_),
    .B1(net203),
    .B2(_12591_),
    .ZN(_12967_));
 OAI21_X2 _22336_ (.A(_12700_),
    .B1(_12948_),
    .B2(_12967_),
    .ZN(_12968_));
 OAI21_X2 _22337_ (.A(_12601_),
    .B1(_12581_),
    .B2(_12676_),
    .ZN(_12969_));
 OAI22_X2 _22338_ (.A1(_12673_),
    .A2(_12851_),
    .B1(_12969_),
    .B2(_12904_),
    .ZN(_12970_));
 OAI33_X1 _22339_ (.A1(_12965_),
    .A2(_12963_),
    .A3(_12968_),
    .B1(_12970_),
    .B2(_12860_),
    .B3(_12638_),
    .ZN(_12971_));
 NAND2_X1 _22340_ (.A1(net140),
    .A2(_12703_),
    .ZN(_12972_));
 OAI21_X1 _22341_ (.A(_12972_),
    .B1(_12652_),
    .B2(net139),
    .ZN(_12973_));
 AND2_X1 _22342_ (.A1(_12842_),
    .A2(_12915_),
    .ZN(_12974_));
 NAND2_X1 _22343_ (.A1(_14956_),
    .A2(_12599_),
    .ZN(_12975_));
 NAND2_X2 _22344_ (.A1(net140),
    .A2(_12550_),
    .ZN(_12976_));
 AND3_X1 _22345_ (.A1(_12691_),
    .A2(_12850_),
    .A3(_12976_),
    .ZN(_12977_));
 AOI221_X2 _22346_ (.A(_12633_),
    .B1(_12973_),
    .B2(_12974_),
    .C1(_12975_),
    .C2(_12977_),
    .ZN(_12978_));
 NAND2_X1 _22347_ (.A1(_12659_),
    .A2(_12881_),
    .ZN(_12979_));
 NOR3_X1 _22348_ (.A1(_12551_),
    .A2(_12796_),
    .A3(_12858_),
    .ZN(_12980_));
 OAI22_X2 _22349_ (.A1(_12856_),
    .A2(_12725_),
    .B1(_12718_),
    .B2(_12546_),
    .ZN(_12981_));
 OAI221_X2 _22350_ (.A(_12757_),
    .B1(_12979_),
    .B2(_12980_),
    .C1(_12981_),
    .C2(_12660_),
    .ZN(_12982_));
 NAND2_X1 _22351_ (.A1(_12722_),
    .A2(_12601_),
    .ZN(_12983_));
 OAI21_X1 _22352_ (.A(_12983_),
    .B1(_12686_),
    .B2(_12695_),
    .ZN(_12984_));
 AOI21_X1 _22353_ (.A(_12638_),
    .B1(_12984_),
    .B2(_12702_),
    .ZN(_12985_));
 AOI221_X2 _22354_ (.A(_12971_),
    .B1(_12978_),
    .B2(_12982_),
    .C1(_12749_),
    .C2(_12985_),
    .ZN(_12986_));
 NOR3_X1 _22355_ (.A1(_14968_),
    .A2(_12654_),
    .A3(_12655_),
    .ZN(_12987_));
 AOI21_X1 _22356_ (.A(_12987_),
    .B1(_12744_),
    .B2(_12701_),
    .ZN(_12988_));
 OAI21_X2 _22357_ (.A(_12567_),
    .B1(_12656_),
    .B2(_12508_),
    .ZN(_12989_));
 OAI22_X2 _22358_ (.A1(_14955_),
    .A2(_12772_),
    .B1(_12966_),
    .B2(_12686_),
    .ZN(_12990_));
 OAI221_X2 _22359_ (.A(_12621_),
    .B1(_12679_),
    .B2(_12988_),
    .C1(_12989_),
    .C2(_12990_),
    .ZN(_12991_));
 OAI221_X1 _22360_ (.A(_12842_),
    .B1(_12703_),
    .B2(_12775_),
    .C1(_14956_),
    .C2(_12708_),
    .ZN(_12992_));
 AOI21_X1 _22361_ (.A(_12547_),
    .B1(_12750_),
    .B2(_12751_),
    .ZN(_12993_));
 NOR3_X1 _22362_ (.A1(_12682_),
    .A2(_12882_),
    .A3(_12724_),
    .ZN(_12994_));
 NAND3_X1 _22363_ (.A1(_12706_),
    .A2(_12691_),
    .A3(_12850_),
    .ZN(_12995_));
 OAI221_X1 _22364_ (.A(_12991_),
    .B1(_12992_),
    .B2(_12993_),
    .C1(_12994_),
    .C2(_12995_),
    .ZN(_12996_));
 OR3_X1 _22365_ (.A1(_12645_),
    .A2(_12719_),
    .A3(_12796_),
    .ZN(_12997_));
 XNOR2_X1 _22366_ (.A(_12775_),
    .B(_12593_),
    .ZN(_12998_));
 OAI211_X2 _22367_ (.A(_12568_),
    .B(_12997_),
    .C1(_12998_),
    .C2(_14972_),
    .ZN(_12999_));
 AOI21_X1 _22368_ (.A(_12679_),
    .B1(_12781_),
    .B2(_14954_),
    .ZN(_13000_));
 AOI21_X1 _22369_ (.A(_12621_),
    .B1(_12851_),
    .B2(_13000_),
    .ZN(_13001_));
 AOI21_X1 _22370_ (.A(_12634_),
    .B1(_12999_),
    .B2(_13001_),
    .ZN(_13002_));
 AND2_X1 _22371_ (.A1(_12701_),
    .A2(_12740_),
    .ZN(_13003_));
 NOR2_X1 _22372_ (.A1(_12724_),
    .A2(_12683_),
    .ZN(_13004_));
 OAI221_X1 _22373_ (.A(_12661_),
    .B1(_13003_),
    .B2(_12969_),
    .C1(_13004_),
    .C2(_12687_),
    .ZN(_13005_));
 OAI21_X1 _22374_ (.A(_12943_),
    .B1(_13003_),
    .B2(_12718_),
    .ZN(_13006_));
 NAND3_X1 _22375_ (.A1(_12622_),
    .A2(_13005_),
    .A3(_13006_),
    .ZN(_13007_));
 AOI22_X1 _22376_ (.A1(_12634_),
    .A2(_12996_),
    .B1(_13002_),
    .B2(_13007_),
    .ZN(_13008_));
 MUX2_X1 _22377_ (.A(_12986_),
    .B(_13008_),
    .S(_12664_),
    .Z(_00076_));
 NAND2_X1 _22378_ (.A1(_12566_),
    .A2(_12608_),
    .ZN(_13009_));
 AOI21_X1 _22379_ (.A(_12606_),
    .B1(_12659_),
    .B2(_12592_),
    .ZN(_13010_));
 AOI221_X2 _22380_ (.A(_12549_),
    .B1(_13009_),
    .B2(_13010_),
    .C1(_12808_),
    .C2(net200),
    .ZN(_13011_));
 AOI22_X2 _22381_ (.A1(net665),
    .A2(_12599_),
    .B1(_12781_),
    .B2(_12549_),
    .ZN(_13012_));
 AOI21_X1 _22382_ (.A(_12781_),
    .B1(_12702_),
    .B2(_12660_),
    .ZN(_13013_));
 OAI221_X2 _22383_ (.A(_12621_),
    .B1(_12661_),
    .B2(_13012_),
    .C1(_13013_),
    .C2(_14960_),
    .ZN(_13014_));
 NAND2_X1 _22384_ (.A1(_12765_),
    .A2(_12846_),
    .ZN(_13015_));
 AOI221_X2 _22385_ (.A(_12567_),
    .B1(_12609_),
    .B2(_12643_),
    .C1(_13015_),
    .C2(_12681_),
    .ZN(_13016_));
 AOI21_X1 _22386_ (.A(_12552_),
    .B1(_12750_),
    .B2(_12762_),
    .ZN(_13017_));
 OAI21_X1 _22387_ (.A(_12679_),
    .B1(_12604_),
    .B2(_14960_),
    .ZN(_13018_));
 OAI21_X1 _22388_ (.A(_12716_),
    .B1(_13017_),
    .B2(_13018_),
    .ZN(_13019_));
 OAI22_X2 _22389_ (.A1(_13011_),
    .A2(_13014_),
    .B1(_13016_),
    .B2(_13019_),
    .ZN(_13020_));
 OAI221_X1 _22390_ (.A(_12757_),
    .B1(_12726_),
    .B2(_12735_),
    .C1(_12708_),
    .C2(_12856_),
    .ZN(_13021_));
 NOR3_X1 _22391_ (.A1(_12667_),
    .A2(_12712_),
    .A3(_13021_),
    .ZN(_13022_));
 AOI22_X2 _22392_ (.A1(_14960_),
    .A2(_12838_),
    .B1(_12786_),
    .B2(_14972_),
    .ZN(_13023_));
 OAI21_X1 _22393_ (.A(_12612_),
    .B1(_13023_),
    .B2(_12622_),
    .ZN(_13024_));
 NOR2_X1 _22394_ (.A1(_14972_),
    .A2(_12715_),
    .ZN(_13025_));
 NOR2_X1 _22395_ (.A1(_12682_),
    .A2(_12715_),
    .ZN(_13026_));
 AOI22_X1 _22396_ (.A1(_12670_),
    .A2(_13025_),
    .B1(_13026_),
    .B2(_12720_),
    .ZN(_13027_));
 AOI21_X1 _22397_ (.A(_13022_),
    .B1(_13024_),
    .B2(_13027_),
    .ZN(_13028_));
 NAND2_X1 _22398_ (.A1(_14979_),
    .A2(_12689_),
    .ZN(_13029_));
 OAI221_X1 _22399_ (.A(_12842_),
    .B1(_12940_),
    .B2(_14979_),
    .C1(_13029_),
    .C2(_14954_),
    .ZN(_13030_));
 NAND2_X1 _22400_ (.A1(_12666_),
    .A2(_13030_),
    .ZN(_13031_));
 OAI221_X1 _22401_ (.A(_12627_),
    .B1(_12666_),
    .B2(_13020_),
    .C1(_13028_),
    .C2(_13031_),
    .ZN(_13032_));
 NAND2_X1 _22402_ (.A1(_12775_),
    .A2(_12725_),
    .ZN(_13033_));
 OAI221_X2 _22403_ (.A(_12667_),
    .B1(_13033_),
    .B2(_12821_),
    .C1(_12933_),
    .C2(_12656_),
    .ZN(_13034_));
 NOR2_X1 _22404_ (.A1(_12735_),
    .A2(_12687_),
    .ZN(_13035_));
 OAI221_X1 _22405_ (.A(_12568_),
    .B1(_12689_),
    .B2(_13035_),
    .C1(_13029_),
    .C2(net138),
    .ZN(_13036_));
 NAND3_X1 _22406_ (.A1(_12622_),
    .A2(_13034_),
    .A3(_13036_),
    .ZN(_13037_));
 OR3_X1 _22407_ (.A1(_12686_),
    .A2(_12684_),
    .A3(_12760_),
    .ZN(_13038_));
 OAI21_X1 _22408_ (.A(_14972_),
    .B1(_12683_),
    .B2(_12797_),
    .ZN(_13039_));
 NAND3_X1 _22409_ (.A1(_12850_),
    .A2(_13038_),
    .A3(_13039_),
    .ZN(_13040_));
 NOR2_X1 _22410_ (.A1(_14979_),
    .A2(_12691_),
    .ZN(_13041_));
 OAI21_X1 _22411_ (.A(_12842_),
    .B1(_13041_),
    .B2(_12684_),
    .ZN(_13042_));
 NAND4_X1 _22412_ (.A1(_12836_),
    .A2(_13037_),
    .A3(_13040_),
    .A4(_13042_),
    .ZN(_13043_));
 OAI33_X1 _22413_ (.A1(_14963_),
    .A2(_12715_),
    .A3(_12882_),
    .B1(_12941_),
    .B2(_12687_),
    .B3(_12676_),
    .ZN(_13044_));
 NAND2_X1 _22414_ (.A1(_12621_),
    .A2(_12726_),
    .ZN(_13045_));
 NAND3_X1 _22415_ (.A1(_14960_),
    .A2(_12715_),
    .A3(_12702_),
    .ZN(_13046_));
 AOI21_X1 _22416_ (.A(_12881_),
    .B1(_13045_),
    .B2(_13046_),
    .ZN(_13047_));
 NOR4_X1 _22417_ (.A1(_12612_),
    .A2(_12756_),
    .A3(_13044_),
    .A4(_13047_),
    .ZN(_13048_));
 NOR2_X1 _22418_ (.A1(_12622_),
    .A2(_12604_),
    .ZN(_13049_));
 OAI21_X1 _22419_ (.A(_14954_),
    .B1(_12599_),
    .B2(_13049_),
    .ZN(_13050_));
 OAI21_X1 _22420_ (.A(_12769_),
    .B1(_12688_),
    .B2(_12775_),
    .ZN(_13051_));
 OR2_X1 _22421_ (.A1(_12686_),
    .A2(_12733_),
    .ZN(_13052_));
 OAI22_X1 _22422_ (.A1(_12682_),
    .A2(_13051_),
    .B1(_13052_),
    .B2(_12904_),
    .ZN(_13053_));
 OR2_X1 _22423_ (.A1(_12688_),
    .A2(_12740_),
    .ZN(_13054_));
 OAI21_X1 _22424_ (.A(_13038_),
    .B1(_13054_),
    .B2(_12682_),
    .ZN(_13055_));
 MUX2_X1 _22425_ (.A(_13053_),
    .B(_13055_),
    .S(_12716_),
    .Z(_13056_));
 NOR2_X1 _22426_ (.A1(_12667_),
    .A2(_12756_),
    .ZN(_13057_));
 AOI22_X1 _22427_ (.A1(_13048_),
    .A2(_13050_),
    .B1(_13056_),
    .B2(_13057_),
    .ZN(_13058_));
 NAND3_X1 _22428_ (.A1(_13032_),
    .A2(_13043_),
    .A3(_13058_),
    .ZN(_00077_));
 NAND2_X1 _22429_ (.A1(_12757_),
    .A2(_12627_),
    .ZN(_13059_));
 NAND2_X1 _22430_ (.A1(_12665_),
    .A2(_12567_),
    .ZN(_13060_));
 AOI21_X1 _22431_ (.A(_13060_),
    .B1(_12599_),
    .B2(_12605_),
    .ZN(_13061_));
 NOR2_X1 _22432_ (.A1(net538),
    .A2(_12701_),
    .ZN(_13062_));
 OAI21_X1 _22433_ (.A(_12552_),
    .B1(_13062_),
    .B2(_12966_),
    .ZN(_13063_));
 NOR2_X1 _22434_ (.A1(net499),
    .A2(_12546_),
    .ZN(_13064_));
 AOI21_X1 _22435_ (.A(_13064_),
    .B1(_12895_),
    .B2(_12645_),
    .ZN(_13065_));
 OAI21_X1 _22436_ (.A(_12897_),
    .B1(_13065_),
    .B2(_12702_),
    .ZN(_13066_));
 AOI221_X2 _22437_ (.A(_13059_),
    .B1(_13061_),
    .B2(_13063_),
    .C1(_12693_),
    .C2(_13066_),
    .ZN(_13067_));
 OR2_X1 _22438_ (.A1(_12552_),
    .A2(_12718_),
    .ZN(_13068_));
 OAI21_X1 _22439_ (.A(_12642_),
    .B1(_12726_),
    .B2(_12775_),
    .ZN(_13069_));
 OAI22_X1 _22440_ (.A1(_12904_),
    .A2(_13068_),
    .B1(_13069_),
    .B2(_12682_),
    .ZN(_13070_));
 NOR3_X1 _22441_ (.A1(_14973_),
    .A2(_14982_),
    .A3(_12688_),
    .ZN(_13071_));
 AOI21_X1 _22442_ (.A(_13071_),
    .B1(_12976_),
    .B2(_12741_),
    .ZN(_13072_));
 MUX2_X1 _22443_ (.A(_13070_),
    .B(_13072_),
    .S(_12666_),
    .Z(_13073_));
 OAI21_X1 _22444_ (.A(_13067_),
    .B1(_13073_),
    .B2(_12612_),
    .ZN(_13074_));
 OAI21_X1 _22445_ (.A(_14972_),
    .B1(_12689_),
    .B2(_12933_),
    .ZN(_13075_));
 OAI221_X1 _22446_ (.A(_12680_),
    .B1(_12831_),
    .B2(_14972_),
    .C1(_13075_),
    .C2(_12904_),
    .ZN(_13076_));
 OAI21_X1 _22447_ (.A(_12689_),
    .B1(_12694_),
    .B2(net200),
    .ZN(_13077_));
 NAND3_X1 _22448_ (.A1(_12650_),
    .A2(_12693_),
    .A3(_13077_),
    .ZN(_13078_));
 NAND4_X1 _22449_ (.A1(_12716_),
    .A2(_12627_),
    .A3(_13076_),
    .A4(_13078_),
    .ZN(_13079_));
 NOR3_X1 _22450_ (.A1(_14979_),
    .A2(_12711_),
    .A3(_12966_),
    .ZN(_13080_));
 NOR2_X1 _22451_ (.A1(_12726_),
    .A2(_12889_),
    .ZN(_13081_));
 NOR3_X1 _22452_ (.A1(_14972_),
    .A2(net911),
    .A3(_13081_),
    .ZN(_13082_));
 OAI21_X1 _22453_ (.A(_12612_),
    .B1(_13080_),
    .B2(_13082_),
    .ZN(_13083_));
 NOR2_X1 _22454_ (.A1(_12605_),
    .A2(_12726_),
    .ZN(_13084_));
 OAI221_X2 _22455_ (.A(_12667_),
    .B1(_13084_),
    .B2(_12962_),
    .C1(_13052_),
    .C2(_13003_),
    .ZN(_13085_));
 AOI21_X1 _22456_ (.A(_12634_),
    .B1(_13083_),
    .B2(_13085_),
    .ZN(_13086_));
 OAI22_X1 _22457_ (.A1(_12676_),
    .A2(_12686_),
    .B1(_12870_),
    .B2(_12695_),
    .ZN(_13087_));
 AOI21_X1 _22458_ (.A(_12679_),
    .B1(_12702_),
    .B2(_13087_),
    .ZN(_13088_));
 MUX2_X1 _22459_ (.A(_12856_),
    .B(net665),
    .S(_12592_),
    .Z(_13089_));
 AOI21_X1 _22460_ (.A(_12989_),
    .B1(_13089_),
    .B2(_12547_),
    .ZN(_13090_));
 NOR2_X1 _22461_ (.A1(_12659_),
    .A2(_12581_),
    .ZN(_13091_));
 AOI211_X2 _22462_ (.A(_12546_),
    .B(_13091_),
    .C1(_12967_),
    .C2(_12659_),
    .ZN(_13092_));
 NAND2_X1 _22463_ (.A1(_12695_),
    .A2(_12567_),
    .ZN(_13093_));
 NAND3_X1 _22464_ (.A1(_12549_),
    .A2(_12860_),
    .A3(_12701_),
    .ZN(_13094_));
 AOI21_X1 _22465_ (.A(_12552_),
    .B1(_13093_),
    .B2(_13094_),
    .ZN(_13095_));
 OAI21_X1 _22466_ (.A(_12665_),
    .B1(_12808_),
    .B2(_14954_),
    .ZN(_13096_));
 OAI33_X1 _22467_ (.A1(_12666_),
    .A2(_13088_),
    .A3(_13090_),
    .B1(_13096_),
    .B2(_13095_),
    .B3(_13092_),
    .ZN(_13097_));
 AOI221_X2 _22468_ (.A(_12566_),
    .B1(_12644_),
    .B2(_12527_),
    .C1(net548),
    .C2(_12505_),
    .ZN(_13098_));
 OAI21_X2 _22469_ (.A(_12791_),
    .B1(_12561_),
    .B2(_12564_),
    .ZN(_13099_));
 OAI33_X1 _22470_ (.A1(_12775_),
    .A2(_12860_),
    .A3(_12703_),
    .B1(_13099_),
    .B2(_12582_),
    .B3(_12644_),
    .ZN(_13100_));
 NOR3_X1 _22471_ (.A1(_12567_),
    .A2(_12725_),
    .A3(_12881_),
    .ZN(_13101_));
 NOR3_X1 _22472_ (.A1(_12549_),
    .A2(_12686_),
    .A3(_12860_),
    .ZN(_13102_));
 NOR4_X1 _22473_ (.A1(_13100_),
    .A2(_13098_),
    .A3(_13101_),
    .A4(_13102_),
    .ZN(_13103_));
 AND2_X1 _22474_ (.A1(_14974_),
    .A2(_12688_),
    .ZN(_13104_));
 NOR2_X1 _22475_ (.A1(_12856_),
    .A2(_12601_),
    .ZN(_13105_));
 AOI211_X2 _22476_ (.A(_12581_),
    .B(_13105_),
    .C1(net723),
    .C2(_12551_),
    .ZN(_13106_));
 OAI21_X1 _22477_ (.A(_12661_),
    .B1(_13104_),
    .B2(_13106_),
    .ZN(_13107_));
 AOI21_X1 _22478_ (.A(_12660_),
    .B1(_12609_),
    .B2(_12643_),
    .ZN(_13108_));
 AOI21_X1 _22479_ (.A(_12665_),
    .B1(_13108_),
    .B2(_12921_),
    .ZN(_13109_));
 AOI22_X1 _22480_ (.A1(_12666_),
    .A2(_13103_),
    .B1(_13107_),
    .B2(_13109_),
    .ZN(_13110_));
 MUX2_X1 _22481_ (.A(_13097_),
    .B(_13110_),
    .S(_12622_),
    .Z(_13111_));
 OAI221_X1 _22482_ (.A(_13074_),
    .B1(_13079_),
    .B2(_13086_),
    .C1(_13111_),
    .C2(_12627_),
    .ZN(_00078_));
 OAI21_X1 _22483_ (.A(net202),
    .B1(_12599_),
    .B2(_12781_),
    .ZN(_13112_));
 AOI22_X1 _22484_ (.A1(_14963_),
    .A2(_12607_),
    .B1(_12609_),
    .B2(net932),
    .ZN(_13113_));
 NAND4_X1 _22485_ (.A1(_12855_),
    .A2(_12850_),
    .A3(_13112_),
    .A4(_13113_),
    .ZN(_13114_));
 NAND2_X1 _22486_ (.A1(_12855_),
    .A2(_12834_),
    .ZN(_13115_));
 OAI21_X1 _22487_ (.A(_12772_),
    .B1(_12751_),
    .B2(_12551_),
    .ZN(_13116_));
 AOI222_X2 _22488_ (.A1(_14956_),
    .A2(_12609_),
    .B1(_13116_),
    .B2(_12775_),
    .C1(_12549_),
    .C2(_12607_),
    .ZN(_13117_));
 NOR2_X1 _22489_ (.A1(_12757_),
    .A2(_12751_),
    .ZN(_13118_));
 NOR3_X1 _22490_ (.A1(_12645_),
    .A2(_12637_),
    .A3(_12760_),
    .ZN(_13119_));
 OAI21_X1 _22491_ (.A(_14960_),
    .B1(_13118_),
    .B2(_13119_),
    .ZN(_13120_));
 NAND3_X1 _22492_ (.A1(_12661_),
    .A2(_12855_),
    .A3(_13120_),
    .ZN(_13121_));
 OAI21_X1 _22493_ (.A(_12856_),
    .B1(_12637_),
    .B2(_12581_),
    .ZN(_13122_));
 MUX2_X1 _22494_ (.A(_12508_),
    .B(_13122_),
    .S(_12828_),
    .Z(_13123_));
 OAI21_X1 _22495_ (.A(_12846_),
    .B1(_12751_),
    .B2(_12620_),
    .ZN(_13124_));
 MUX2_X1 _22496_ (.A(_13123_),
    .B(_13124_),
    .S(_12552_),
    .Z(_13125_));
 OAI221_X2 _22497_ (.A(_13114_),
    .B1(_13115_),
    .B2(_13117_),
    .C1(_13121_),
    .C2(_13125_),
    .ZN(_13126_));
 NOR2_X1 _22498_ (.A1(_12527_),
    .A2(_13009_),
    .ZN(_13127_));
 AOI21_X1 _22499_ (.A(_12607_),
    .B1(_12581_),
    .B2(_12658_),
    .ZN(_13128_));
 NOR2_X1 _22500_ (.A1(_12549_),
    .A2(_13128_),
    .ZN(_13129_));
 OAI21_X1 _22501_ (.A(_12775_),
    .B1(_13127_),
    .B2(_13129_),
    .ZN(_13130_));
 AOI221_X2 _22502_ (.A(_12620_),
    .B1(_12658_),
    .B2(_12545_),
    .C1(_12781_),
    .C2(net203),
    .ZN(_13131_));
 NOR2_X1 _22503_ (.A1(net139),
    .A2(_12772_),
    .ZN(_13132_));
 AOI21_X1 _22504_ (.A(net722),
    .B1(_12708_),
    .B2(_12751_),
    .ZN(_13133_));
 OAI21_X1 _22505_ (.A(_12860_),
    .B1(_13132_),
    .B2(_13133_),
    .ZN(_13134_));
 AOI21_X1 _22506_ (.A(_12668_),
    .B1(_12608_),
    .B2(_12549_),
    .ZN(_13135_));
 AOI21_X1 _22507_ (.A(_12599_),
    .B1(_12781_),
    .B2(_12527_),
    .ZN(_13136_));
 OAI221_X2 _22508_ (.A(_13134_),
    .B1(_13135_),
    .B2(_12860_),
    .C1(_12695_),
    .C2(_13136_),
    .ZN(_13137_));
 AOI221_X2 _22509_ (.A(_12819_),
    .B1(_13130_),
    .B2(_13131_),
    .C1(_13137_),
    .C2(_12757_),
    .ZN(_13138_));
 NOR2_X1 _22510_ (.A1(_12622_),
    .A2(_12666_),
    .ZN(_13139_));
 OR2_X1 _22511_ (.A1(_14982_),
    .A2(_12593_),
    .ZN(_13140_));
 NAND2_X1 _22512_ (.A1(_12705_),
    .A2(_12686_),
    .ZN(_13141_));
 NAND3_X1 _22513_ (.A1(_12726_),
    .A2(_12646_),
    .A3(_13141_),
    .ZN(_13142_));
 NAND3_X1 _22514_ (.A1(_12661_),
    .A2(_13140_),
    .A3(_13142_),
    .ZN(_13143_));
 OAI21_X1 _22515_ (.A(_12769_),
    .B1(_12688_),
    .B2(net200),
    .ZN(_13144_));
 AOI21_X1 _22516_ (.A(_12764_),
    .B1(_13144_),
    .B2(_12687_),
    .ZN(_13145_));
 OAI21_X1 _22517_ (.A(_13143_),
    .B1(_13145_),
    .B2(_12667_),
    .ZN(_13146_));
 AOI21_X2 _22518_ (.A(_12664_),
    .B1(_13139_),
    .B2(_13146_),
    .ZN(_13147_));
 MUX2_X1 _22519_ (.A(_12676_),
    .B(net723),
    .S(_12546_),
    .Z(_13148_));
 OAI221_X1 _22520_ (.A(_12679_),
    .B1(_13033_),
    .B2(_12694_),
    .C1(_13148_),
    .C2(_12726_),
    .ZN(_13149_));
 NAND2_X1 _22521_ (.A1(_12605_),
    .A2(_12645_),
    .ZN(_13150_));
 MUX2_X1 _22522_ (.A(_14968_),
    .B(_13150_),
    .S(_12593_),
    .Z(_13151_));
 OAI21_X1 _22523_ (.A(_13149_),
    .B1(_13151_),
    .B2(_12568_),
    .ZN(_13152_));
 AOI22_X1 _22524_ (.A1(_12735_),
    .A2(_12593_),
    .B1(_12741_),
    .B2(_12976_),
    .ZN(_13153_));
 OR2_X1 _22525_ (.A1(_12845_),
    .A2(_13153_),
    .ZN(_13154_));
 NOR2_X1 _22526_ (.A1(_12601_),
    .A2(_12684_),
    .ZN(_13155_));
 AOI221_X2 _22527_ (.A(_12837_),
    .B1(_13155_),
    .B2(_12691_),
    .C1(_12551_),
    .C2(_12798_),
    .ZN(_13156_));
 NAND3_X1 _22528_ (.A1(_12637_),
    .A2(_12659_),
    .A3(_12983_),
    .ZN(_13157_));
 AOI21_X1 _22529_ (.A(_13157_),
    .B1(_12759_),
    .B2(_12820_),
    .ZN(_13158_));
 AOI22_X1 _22530_ (.A1(net547),
    .A2(_12505_),
    .B1(_12548_),
    .B2(_12545_),
    .ZN(_13159_));
 OAI221_X1 _22531_ (.A(_12620_),
    .B1(_12561_),
    .B2(_12564_),
    .C1(_12582_),
    .C2(_13159_),
    .ZN(_13160_));
 AOI21_X1 _22532_ (.A(_13160_),
    .B1(_12934_),
    .B2(_12688_),
    .ZN(_13161_));
 NOR4_X2 _22533_ (.A1(_13161_),
    .A2(_12634_),
    .A3(_13158_),
    .A4(_13156_),
    .ZN(_13162_));
 AOI22_X2 _22534_ (.A1(_12700_),
    .A2(_13152_),
    .B1(_13162_),
    .B2(_13154_),
    .ZN(_13163_));
 AOI211_X2 _22535_ (.A(_13126_),
    .B(_13138_),
    .C1(_13163_),
    .C2(_13147_),
    .ZN(_00079_));
 INV_X1 _22536_ (.A(_06260_),
    .ZN(_13164_));
 NOR2_X1 _22537_ (.A1(_13164_),
    .A2(_08995_),
    .ZN(_13165_));
 NOR2_X1 _22538_ (.A1(_06260_),
    .A2(_08995_),
    .ZN(_13166_));
 XNOR2_X2 _22539_ (.A(\sa02_sr[1] ),
    .B(\sa31_sub[1] ),
    .ZN(_13167_));
 XNOR2_X2 _22540_ (.A(_13167_),
    .B(_10504_),
    .ZN(_13168_));
 XNOR2_X2 _22541_ (.A(_10455_),
    .B(\sa20_sub[1] ),
    .ZN(_13169_));
 XNOR2_X2 _22542_ (.A(_13169_),
    .B(_13168_),
    .ZN(_13170_));
 MUX2_X2 _22543_ (.A(_13165_),
    .B(_13166_),
    .S(_13170_),
    .Z(_13171_));
 NAND3_X4 _22544_ (.A1(_06260_),
    .A2(_09818_),
    .A3(_00458_),
    .ZN(_13172_));
 NAND2_X4 _22545_ (.A1(_09818_),
    .A2(_13164_),
    .ZN(_13173_));
 OAI21_X4 _22546_ (.A(_13172_),
    .B1(_00458_),
    .B2(_13173_),
    .ZN(_13174_));
 NOR2_X4 _22547_ (.A1(_13174_),
    .A2(_13171_),
    .ZN(_13175_));
 INV_X8 _22548_ (.A(net487),
    .ZN(_13176_));
 BUF_X16 _22549_ (.A(_13176_),
    .Z(_13177_));
 BUF_X16 _22550_ (.A(_13177_),
    .Z(_13178_));
 BUF_X16 _22551_ (.A(_13178_),
    .Z(_14992_));
 XNOR2_X2 _22552_ (.A(_10439_),
    .B(_10453_),
    .ZN(_13179_));
 XNOR2_X1 _22553_ (.A(net621),
    .B(_13179_),
    .ZN(_13180_));
 XOR2_X2 _22554_ (.A(net550),
    .B(_10503_),
    .Z(_13181_));
 NAND3_X1 _22555_ (.A1(_06247_),
    .A2(_09074_),
    .A3(_13181_),
    .ZN(_13182_));
 NOR2_X1 _22556_ (.A1(_06247_),
    .A2(_08972_),
    .ZN(_13183_));
 NAND2_X1 _22557_ (.A1(net521),
    .A2(_13183_),
    .ZN(_13184_));
 AOI21_X1 _22558_ (.A(_13180_),
    .B1(_13182_),
    .B2(_13184_),
    .ZN(_13185_));
 XOR2_X2 _22559_ (.A(_10439_),
    .B(_10453_),
    .Z(_13186_));
 XNOR2_X1 _22560_ (.A(net597),
    .B(_13186_),
    .ZN(_13187_));
 NAND2_X1 _22561_ (.A1(_13181_),
    .A2(_13183_),
    .ZN(_13188_));
 NAND3_X1 _22562_ (.A1(_06247_),
    .A2(_09099_),
    .A3(net521),
    .ZN(_13189_));
 AOI21_X1 _22563_ (.A(_13187_),
    .B1(_13188_),
    .B2(_13189_),
    .ZN(_13190_));
 INV_X1 _22564_ (.A(_06247_),
    .ZN(_13191_));
 NAND3_X1 _22565_ (.A1(_13191_),
    .A2(_09015_),
    .A3(_00459_),
    .ZN(_13192_));
 NAND2_X1 _22566_ (.A1(_06247_),
    .A2(_08993_),
    .ZN(_13193_));
 OAI21_X1 _22567_ (.A(_13192_),
    .B1(_13193_),
    .B2(_00459_),
    .ZN(_13194_));
 OR3_X1 _22568_ (.A1(_13185_),
    .A2(_13190_),
    .A3(_13194_),
    .ZN(_13195_));
 BUF_X4 _22569_ (.A(_13195_),
    .Z(_13196_));
 INV_X4 _22570_ (.A(_13196_),
    .ZN(_13197_));
 BUF_X4 _22571_ (.A(_13197_),
    .Z(_14995_));
 XNOR2_X2 _22572_ (.A(_10475_),
    .B(_10550_),
    .ZN(_13198_));
 XNOR2_X1 _22573_ (.A(_10479_),
    .B(_13198_),
    .ZN(_13199_));
 XOR2_X2 _22574_ (.A(net532),
    .B(net557),
    .Z(_13200_));
 NAND3_X1 _22575_ (.A1(_06299_),
    .A2(_09009_),
    .A3(_13200_),
    .ZN(_13201_));
 NOR2_X1 _22576_ (.A1(_06299_),
    .A2(_08970_),
    .ZN(_13202_));
 NAND2_X1 _22577_ (.A1(net711),
    .A2(_13202_),
    .ZN(_13203_));
 AOI21_X2 _22578_ (.A(_13199_),
    .B1(_13201_),
    .B2(_13203_),
    .ZN(_13204_));
 XOR2_X2 _22579_ (.A(_10475_),
    .B(_10550_),
    .Z(_13205_));
 XNOR2_X1 _22580_ (.A(_10479_),
    .B(_13205_),
    .ZN(_13206_));
 NAND2_X1 _22581_ (.A1(_13200_),
    .A2(_13202_),
    .ZN(_13207_));
 NAND3_X1 _22582_ (.A1(_06299_),
    .A2(_09009_),
    .A3(net711),
    .ZN(_13208_));
 AOI21_X2 _22583_ (.A(_13206_),
    .B1(_13207_),
    .B2(_13208_),
    .ZN(_13209_));
 NAND3_X1 _22584_ (.A1(_06306_),
    .A2(net587),
    .A3(_00460_),
    .ZN(_13210_));
 NAND2_X1 _22585_ (.A1(_06299_),
    .A2(net587),
    .ZN(_13211_));
 OAI21_X2 _22586_ (.A(_13210_),
    .B1(_13211_),
    .B2(_00460_),
    .ZN(_13212_));
 NOR3_X4 _22587_ (.A1(_13204_),
    .A2(_13209_),
    .A3(_13212_),
    .ZN(_13213_));
 INV_X2 _22588_ (.A(_13213_),
    .ZN(_13214_));
 BUF_X4 _22589_ (.A(_13214_),
    .Z(_13215_));
 BUF_X4 _22590_ (.A(_13215_),
    .Z(_13216_));
 BUF_X4 _22591_ (.A(_13216_),
    .Z(_13217_));
 CLKBUF_X3 _22592_ (.A(_13217_),
    .Z(_13218_));
 BUF_X4 _22593_ (.A(_13218_),
    .Z(_15011_));
 BUF_X4 _22594_ (.A(_13196_),
    .Z(_13219_));
 BUF_X4 _22595_ (.A(_13219_),
    .Z(_14986_));
 BUF_X4 _22596_ (.A(_13213_),
    .Z(_13220_));
 BUF_X4 _22597_ (.A(_13220_),
    .Z(_13221_));
 BUF_X4 _22598_ (.A(_13221_),
    .Z(_13222_));
 BUF_X4 _22599_ (.A(_13222_),
    .Z(_13223_));
 BUF_X4 _22600_ (.A(_13223_),
    .Z(_15004_));
 XNOR2_X2 _22601_ (.A(_10432_),
    .B(_10506_),
    .ZN(_13224_));
 XNOR2_X1 _22602_ (.A(_10514_),
    .B(net710),
    .ZN(_13225_));
 XNOR2_X1 _22603_ (.A(_10503_),
    .B(_13225_),
    .ZN(_13226_));
 MUX2_X2 _22604_ (.A(\text_in_r[55] ),
    .B(_13226_),
    .S(_09175_),
    .Z(_13227_));
 XNOR2_X2 _22605_ (.A(_06590_),
    .B(_13227_),
    .ZN(_13228_));
 XNOR2_X2 _22606_ (.A(_10512_),
    .B(_10505_),
    .ZN(_13229_));
 XNOR2_X1 _22607_ (.A(_10523_),
    .B(_10513_),
    .ZN(_13230_));
 XNOR2_X1 _22608_ (.A(_13229_),
    .B(_13230_),
    .ZN(_13231_));
 XNOR2_X1 _22609_ (.A(_10515_),
    .B(_13231_),
    .ZN(_13232_));
 MUX2_X2 _22610_ (.A(\text_in_r[54] ),
    .B(_13232_),
    .S(_11191_),
    .Z(_13233_));
 XOR2_X2 _22611_ (.A(_06578_),
    .B(_13233_),
    .Z(_13234_));
 BUF_X4 _22612_ (.A(_13234_),
    .Z(_13235_));
 NOR2_X2 _22613_ (.A1(_13228_),
    .A2(_13235_),
    .ZN(_13236_));
 BUF_X4 _22614_ (.A(_13216_),
    .Z(_13237_));
 CLKBUF_X3 _22615_ (.A(_13237_),
    .Z(_13238_));
 BUF_X4 clone141 (.A(net1),
    .Z(net141));
 BUF_X4 _22617_ (.A(_14990_),
    .Z(_13240_));
 NAND2_X1 _22618_ (.A1(_06228_),
    .A2(net947),
    .ZN(_13241_));
 INV_X1 _22619_ (.A(_06228_),
    .ZN(_13242_));
 NAND2_X1 _22620_ (.A1(_13242_),
    .A2(net947),
    .ZN(_13243_));
 XNOR2_X1 _22621_ (.A(_10480_),
    .B(net522),
    .ZN(_13244_));
 XOR2_X1 _22622_ (.A(_10554_),
    .B(_10535_),
    .Z(_13245_));
 XNOR2_X1 _22623_ (.A(_10551_),
    .B(_13245_),
    .ZN(_13246_));
 XNOR2_X1 _22624_ (.A(_13244_),
    .B(_13246_),
    .ZN(_13247_));
 MUX2_X1 _22625_ (.A(_13241_),
    .B(_13243_),
    .S(_13247_),
    .Z(_13248_));
 BUF_X8 _22626_ (.A(_13248_),
    .Z(_13249_));
 OR3_X2 _22627_ (.A1(_13242_),
    .A2(net948),
    .A3(\text_in_r[51] ),
    .ZN(_13250_));
 NAND3_X2 _22628_ (.A1(_13242_),
    .A2(_09027_),
    .A3(\text_in_r[51] ),
    .ZN(_13251_));
 AND2_X1 _22629_ (.A1(_13250_),
    .A2(_13251_),
    .ZN(_13252_));
 BUF_X8 _22630_ (.A(_13252_),
    .Z(_13253_));
 NAND2_X1 _22631_ (.A1(_13249_),
    .A2(_13253_),
    .ZN(_13254_));
 BUF_X4 _22632_ (.A(_13254_),
    .Z(_13255_));
 BUF_X8 _22633_ (.A(_13255_),
    .Z(_13256_));
 BUF_X4 _22634_ (.A(_13256_),
    .Z(_13257_));
 NOR2_X1 _22635_ (.A1(_13240_),
    .A2(_13257_),
    .ZN(_13258_));
 NOR2_X1 _22636_ (.A1(_13242_),
    .A2(_09726_),
    .ZN(_13259_));
 NOR2_X1 _22637_ (.A1(_06228_),
    .A2(_09726_),
    .ZN(_13260_));
 MUX2_X2 _22638_ (.A(_13259_),
    .B(_13260_),
    .S(_13247_),
    .Z(_13261_));
 BUF_X8 _22639_ (.A(_13261_),
    .Z(_13262_));
 NAND2_X4 _22640_ (.A1(_13250_),
    .A2(_13251_),
    .ZN(_13263_));
 OAI21_X4 _22641_ (.A(_13196_),
    .B1(_13262_),
    .B2(_13263_),
    .ZN(_13264_));
 NOR2_X2 _22642_ (.A1(net174),
    .A2(_13264_),
    .ZN(_13265_));
 NOR3_X1 _22643_ (.A1(_13238_),
    .A2(_13258_),
    .A3(_13265_),
    .ZN(_13266_));
 XNOR2_X1 _22644_ (.A(_10541_),
    .B(_10503_),
    .ZN(_13267_));
 XNOR2_X1 _22645_ (.A(_10551_),
    .B(_13267_),
    .ZN(_13268_));
 XOR2_X1 _22646_ (.A(_10536_),
    .B(_10527_),
    .Z(_13269_));
 XNOR2_X1 _22647_ (.A(_10540_),
    .B(_13269_),
    .ZN(_13270_));
 XNOR2_X1 _22648_ (.A(_13268_),
    .B(_13270_),
    .ZN(_13271_));
 MUX2_X2 _22649_ (.A(\text_in_r[52] ),
    .B(_13271_),
    .S(_09023_),
    .Z(_13272_));
 XNOR2_X2 _22650_ (.A(_06284_),
    .B(_13272_),
    .ZN(_13273_));
 BUF_X4 _22651_ (.A(_13273_),
    .Z(_13274_));
 BUF_X4 _22652_ (.A(_13274_),
    .Z(_13275_));
 BUF_X4 _22653_ (.A(_13275_),
    .Z(_13276_));
 BUF_X4 _22654_ (.A(_14998_),
    .Z(_13277_));
 AOI21_X4 _22655_ (.A(_13213_),
    .B1(_13249_),
    .B2(_13253_),
    .ZN(_13278_));
 NAND2_X1 _22656_ (.A1(_13277_),
    .A2(_13278_),
    .ZN(_13279_));
 NAND2_X1 _22657_ (.A1(_13276_),
    .A2(_13279_),
    .ZN(_13280_));
 NOR2_X4 _22658_ (.A1(_13262_),
    .A2(_13263_),
    .ZN(_13281_));
 BUF_X4 _22659_ (.A(_13281_),
    .Z(_13282_));
 NAND3_X4 _22660_ (.A1(_13196_),
    .A2(_13249_),
    .A3(_13253_),
    .ZN(_13283_));
 BUF_X8 _22661_ (.A(_13175_),
    .Z(_13284_));
 OAI221_X2 _22662_ (.A(_13222_),
    .B1(_13282_),
    .B2(_13240_),
    .C1(_13283_),
    .C2(net1),
    .ZN(_13285_));
 BUF_X4 _22663_ (.A(_13249_),
    .Z(_13286_));
 BUF_X4 _22664_ (.A(_13253_),
    .Z(_13287_));
 NAND3_X4 _22665_ (.A1(_13214_),
    .A2(_13286_),
    .A3(_13287_),
    .ZN(_13288_));
 BUF_X4 _22666_ (.A(_14996_),
    .Z(_13289_));
 OAI21_X1 _22667_ (.A(_13285_),
    .B1(_13288_),
    .B2(_13289_),
    .ZN(_13290_));
 OAI221_X1 _22668_ (.A(_13236_),
    .B1(_13266_),
    .B2(_13280_),
    .C1(_13290_),
    .C2(_13276_),
    .ZN(_13291_));
 XNOR2_X1 _22669_ (.A(_10536_),
    .B(_10516_),
    .ZN(_13292_));
 XNOR2_X1 _22670_ (.A(_10525_),
    .B(_13292_),
    .ZN(_13293_));
 XNOR2_X1 _22671_ (.A(_10526_),
    .B(_13293_),
    .ZN(_13294_));
 MUX2_X2 _22672_ (.A(\text_in_r[53] ),
    .B(_13294_),
    .S(net947),
    .Z(_13295_));
 XNOR2_X2 _22673_ (.A(_06272_),
    .B(_13295_),
    .ZN(_13296_));
 BUF_X4 _22674_ (.A(_13296_),
    .Z(_13297_));
 BUF_X4 _22675_ (.A(_13297_),
    .Z(_13298_));
 XOR2_X2 _22676_ (.A(_06284_),
    .B(_13272_),
    .Z(_13299_));
 BUF_X4 _22677_ (.A(_13299_),
    .Z(_13300_));
 XOR2_X2 _22678_ (.A(_06590_),
    .B(_13227_),
    .Z(_13301_));
 NAND2_X2 _22679_ (.A1(_13301_),
    .A2(_13234_),
    .ZN(_13302_));
 NOR2_X1 _22680_ (.A1(_13300_),
    .A2(_13302_),
    .ZN(_13303_));
 AOI21_X2 _22681_ (.A(_13289_),
    .B1(_13286_),
    .B2(_13287_),
    .ZN(_13304_));
 BUF_X4 _22682_ (.A(_14989_),
    .Z(_13305_));
 NOR3_X4 _22683_ (.A1(_13305_),
    .A2(_13262_),
    .A3(_13263_),
    .ZN(_13306_));
 NOR3_X1 _22684_ (.A1(_13221_),
    .A2(_13304_),
    .A3(_13306_),
    .ZN(_13307_));
 MUX2_X1 _22685_ (.A(net173),
    .B(_13219_),
    .S(_13255_),
    .Z(_13308_));
 BUF_X4 _22686_ (.A(_13220_),
    .Z(_13309_));
 AOI21_X1 _22687_ (.A(_13307_),
    .B1(_13308_),
    .B2(_13309_),
    .ZN(_13310_));
 NAND3_X2 _22688_ (.A1(_14990_),
    .A2(_13249_),
    .A3(_13253_),
    .ZN(_13311_));
 BUF_X2 clone143 (.A(_15125_),
    .Z(net143));
 OAI21_X4 _22690_ (.A(net489),
    .B1(_13262_),
    .B2(_13263_),
    .ZN(_13313_));
 AND3_X4 _22691_ (.A1(_13220_),
    .A2(_13311_),
    .A3(_13313_),
    .ZN(_13314_));
 BUF_X8 _22692_ (.A(_13262_),
    .Z(_13315_));
 BUF_X8 _22693_ (.A(_13263_),
    .Z(_13316_));
 NOR3_X4 _22694_ (.A1(_13220_),
    .A2(_13315_),
    .A3(_13316_),
    .ZN(_13317_));
 CLKBUF_X2 split189 (.A(net896),
    .Z(net189));
 AOI21_X2 _22696_ (.A(_13314_),
    .B1(_13317_),
    .B2(_14988_),
    .ZN(_13319_));
 NOR2_X1 _22697_ (.A1(_13275_),
    .A2(_13302_),
    .ZN(_13320_));
 AOI221_X2 _22698_ (.A(_13298_),
    .B1(_13303_),
    .B2(_13310_),
    .C1(_13319_),
    .C2(_13320_),
    .ZN(_13321_));
 AND2_X1 _22699_ (.A1(_13291_),
    .A2(_13321_),
    .ZN(_13322_));
 XNOR2_X2 _22700_ (.A(_06578_),
    .B(_13233_),
    .ZN(_13323_));
 NOR2_X2 _22701_ (.A1(_13323_),
    .A2(_13300_),
    .ZN(_13324_));
 NOR2_X2 _22702_ (.A1(_13176_),
    .A2(_13281_),
    .ZN(_13325_));
 NAND2_X1 _22703_ (.A1(_14986_),
    .A2(_13218_),
    .ZN(_13326_));
 OAI21_X2 _22704_ (.A(_13220_),
    .B1(_13315_),
    .B2(_13316_),
    .ZN(_13327_));
 BUF_X4 _22705_ (.A(_13327_),
    .Z(_13328_));
 BUF_X8 _22706_ (.A(_14993_),
    .Z(_13329_));
 OAI22_X1 _22707_ (.A1(_13325_),
    .A2(_13326_),
    .B1(_13328_),
    .B2(net540),
    .ZN(_13330_));
 AOI21_X1 _22708_ (.A(_13301_),
    .B1(_13324_),
    .B2(_13330_),
    .ZN(_13331_));
 INV_X8 _22709_ (.A(_13305_),
    .ZN(_13332_));
 NAND3_X2 _22710_ (.A1(_13332_),
    .A2(_13249_),
    .A3(_13253_),
    .ZN(_13333_));
 CLKBUF_X3 _22711_ (.A(_13256_),
    .Z(_13334_));
 NAND2_X1 _22712_ (.A1(_13289_),
    .A2(_13334_),
    .ZN(_13335_));
 AOI21_X1 _22713_ (.A(_13238_),
    .B1(_13333_),
    .B2(_13335_),
    .ZN(_13336_));
 CLKBUF_X3 _22714_ (.A(_13309_),
    .Z(_13337_));
 CLKBUF_X3 _22715_ (.A(_13337_),
    .Z(_13338_));
 NOR3_X4 _22716_ (.A1(_13219_),
    .A2(_13315_),
    .A3(_13316_),
    .ZN(_13339_));
 NAND2_X2 _22717_ (.A1(_13178_),
    .A2(_13339_),
    .ZN(_13340_));
 NAND2_X1 _22718_ (.A1(_14988_),
    .A2(_13334_),
    .ZN(_13341_));
 AOI21_X1 _22719_ (.A(_13338_),
    .B1(_13340_),
    .B2(_13341_),
    .ZN(_13342_));
 NOR2_X1 _22720_ (.A1(_13336_),
    .A2(_13342_),
    .ZN(_13343_));
 NAND2_X2 _22721_ (.A1(_13323_),
    .A2(_13275_),
    .ZN(_13344_));
 BUF_X4 _22722_ (.A(_13276_),
    .Z(_13345_));
 BUF_X4 _22723_ (.A(_13282_),
    .Z(_13346_));
 CLKBUF_X3 _22724_ (.A(_13346_),
    .Z(_13347_));
 CLKBUF_X3 _22725_ (.A(_13309_),
    .Z(_13348_));
 AOI21_X1 _22726_ (.A(_14986_),
    .B1(_13348_),
    .B2(_13323_),
    .ZN(_13349_));
 OAI21_X2 _22727_ (.A(_13219_),
    .B1(_13174_),
    .B2(_13171_),
    .ZN(_13350_));
 NOR2_X1 _22728_ (.A1(_13235_),
    .A2(_13350_),
    .ZN(_13351_));
 OAI21_X1 _22729_ (.A(_13347_),
    .B1(_13349_),
    .B2(_13351_),
    .ZN(_13352_));
 BUF_X4 _22730_ (.A(_13305_),
    .Z(_13353_));
 MUX2_X1 _22731_ (.A(_13353_),
    .B(_14995_),
    .S(_13323_),
    .Z(_13354_));
 BUF_X4 _22732_ (.A(_15002_),
    .Z(_13355_));
 INV_X8 _22733_ (.A(_13355_),
    .ZN(_13356_));
 NOR2_X2 _22734_ (.A1(_13356_),
    .A2(_13221_),
    .ZN(_13357_));
 AOI22_X2 _22735_ (.A1(_13223_),
    .A2(_13354_),
    .B1(_13357_),
    .B2(_13235_),
    .ZN(_13358_));
 MUX2_X1 _22736_ (.A(_13264_),
    .B(_13288_),
    .S(_13235_),
    .Z(_13359_));
 OAI221_X2 _22737_ (.A(_13352_),
    .B1(_13358_),
    .B2(_13347_),
    .C1(net178),
    .C2(_13359_),
    .ZN(_13360_));
 OAI221_X2 _22738_ (.A(_13331_),
    .B1(_13343_),
    .B2(_13344_),
    .C1(_13345_),
    .C2(_13360_),
    .ZN(_13361_));
 BUF_X4 _22739_ (.A(_13300_),
    .Z(_13362_));
 BUF_X4 _22740_ (.A(_13362_),
    .Z(_13363_));
 BUF_X4 _22741_ (.A(_13235_),
    .Z(_13364_));
 NOR2_X1 _22742_ (.A1(_13356_),
    .A2(_13346_),
    .ZN(_13365_));
 NOR2_X2 _22743_ (.A1(_13175_),
    .A2(_13255_),
    .ZN(_13366_));
 NOR3_X1 _22744_ (.A1(_13238_),
    .A2(_13365_),
    .A3(_13366_),
    .ZN(_13367_));
 NOR2_X4 _22745_ (.A1(_13176_),
    .A2(_13255_),
    .ZN(_13368_));
 NOR2_X1 _22746_ (.A1(_13368_),
    .A2(_13326_),
    .ZN(_13369_));
 OAI21_X1 _22747_ (.A(_13364_),
    .B1(_13367_),
    .B2(_13369_),
    .ZN(_13370_));
 BUF_X4 _22748_ (.A(_13323_),
    .Z(_13371_));
 NAND3_X4 _22749_ (.A1(_13305_),
    .A2(_13249_),
    .A3(_13253_),
    .ZN(_13372_));
 NOR2_X1 _22750_ (.A1(net178),
    .A2(_13223_),
    .ZN(_13373_));
 NAND2_X1 _22751_ (.A1(net611),
    .A2(_13238_),
    .ZN(_13374_));
 OAI221_X1 _22752_ (.A(_13371_),
    .B1(_13372_),
    .B2(_13373_),
    .C1(_13374_),
    .C2(_13368_),
    .ZN(_13375_));
 NAND3_X1 _22753_ (.A1(_13363_),
    .A2(_13370_),
    .A3(_13375_),
    .ZN(_13376_));
 XOR2_X2 _22754_ (.A(_06272_),
    .B(_13295_),
    .Z(_13377_));
 BUF_X4 _22755_ (.A(_13377_),
    .Z(_13378_));
 BUF_X4 _22756_ (.A(_13378_),
    .Z(_13379_));
 NOR2_X1 _22757_ (.A1(_13289_),
    .A2(_13288_),
    .ZN(_13380_));
 AOI21_X4 _22758_ (.A(_13215_),
    .B1(_13286_),
    .B2(_13287_),
    .ZN(_13381_));
 OAI21_X4 _22759_ (.A(_13215_),
    .B1(_13315_),
    .B2(_13316_),
    .ZN(_13382_));
 NAND3_X4 _22760_ (.A1(_13213_),
    .A2(_13249_),
    .A3(_13253_),
    .ZN(_13383_));
 NAND2_X2 _22761_ (.A1(_13382_),
    .A2(_13383_),
    .ZN(_13384_));
 INV_X2 _22762_ (.A(_14988_),
    .ZN(_13385_));
 AOI221_X2 _22763_ (.A(_13380_),
    .B1(_13381_),
    .B2(net612),
    .C1(_13384_),
    .C2(_13385_),
    .ZN(_13386_));
 OAI221_X1 _22764_ (.A(_13324_),
    .B1(_13383_),
    .B2(_13240_),
    .C1(_14995_),
    .C2(_13382_),
    .ZN(_13387_));
 BUF_X1 rebuffer138 (.A(_09002_),
    .Z(net632));
 AOI21_X1 _22766_ (.A(_13317_),
    .B1(_13381_),
    .B2(_14995_),
    .ZN(_13389_));
 NOR2_X1 _22767_ (.A1(_13284_),
    .A2(_13389_),
    .ZN(_13390_));
 OAI22_X1 _22768_ (.A1(_13344_),
    .A2(_13386_),
    .B1(_13387_),
    .B2(_13390_),
    .ZN(_13391_));
 NOR3_X1 _22769_ (.A1(_13301_),
    .A2(_13379_),
    .A3(_13391_),
    .ZN(_13392_));
 CLKBUF_X3 _22770_ (.A(_13257_),
    .Z(_13393_));
 AOI22_X1 _22771_ (.A1(_15009_),
    .A2(_13393_),
    .B1(_13317_),
    .B2(_13353_),
    .ZN(_13394_));
 AOI21_X1 _22772_ (.A(_13364_),
    .B1(_13363_),
    .B2(_13394_),
    .ZN(_13395_));
 NAND2_X2 _22773_ (.A1(_13219_),
    .A2(_13220_),
    .ZN(_13396_));
 OAI22_X4 _22774_ (.A1(_13329_),
    .A2(_13309_),
    .B1(_13396_),
    .B2(net1),
    .ZN(_13397_));
 OAI21_X2 _22775_ (.A(_13275_),
    .B1(_13334_),
    .B2(_13397_),
    .ZN(_13398_));
 OAI21_X4 _22776_ (.A(_13197_),
    .B1(_13315_),
    .B2(_13316_),
    .ZN(_13399_));
 NAND2_X1 _22777_ (.A1(_13311_),
    .A2(_13399_),
    .ZN(_13400_));
 NAND2_X1 _22778_ (.A1(_13238_),
    .A2(_13400_),
    .ZN(_13401_));
 OAI21_X1 _22779_ (.A(_13401_),
    .B1(_13328_),
    .B2(_14988_),
    .ZN(_13402_));
 OAI21_X1 _22780_ (.A(_13395_),
    .B1(_13398_),
    .B2(_13402_),
    .ZN(_13403_));
 NAND2_X2 _22781_ (.A1(_13301_),
    .A2(_13297_),
    .ZN(_13404_));
 NOR2_X2 _22782_ (.A1(net612),
    .A2(_13282_),
    .ZN(_13405_));
 NOR3_X4 _22783_ (.A1(_13277_),
    .A2(_13315_),
    .A3(_13316_),
    .ZN(_13406_));
 OAI21_X1 _22784_ (.A(_13337_),
    .B1(_13405_),
    .B2(_13406_),
    .ZN(_13407_));
 NAND2_X1 _22785_ (.A1(_13234_),
    .A2(_13300_),
    .ZN(_13408_));
 NOR2_X2 _22786_ (.A1(_13329_),
    .A2(_13288_),
    .ZN(_13409_));
 NOR2_X1 _22787_ (.A1(_13408_),
    .A2(_13409_),
    .ZN(_13410_));
 INV_X1 _22788_ (.A(_13174_),
    .ZN(_13411_));
 NAND2_X1 _22789_ (.A1(_06260_),
    .A2(_10571_),
    .ZN(_13412_));
 NAND2_X1 _22790_ (.A1(_13164_),
    .A2(_10571_),
    .ZN(_13413_));
 MUX2_X2 _22791_ (.A(_13412_),
    .B(_13413_),
    .S(_13170_),
    .Z(_13414_));
 AOI21_X4 _22792_ (.A(_13196_),
    .B1(_13411_),
    .B2(_13414_),
    .ZN(_13415_));
 NOR2_X1 _22793_ (.A1(_13282_),
    .A2(_13415_),
    .ZN(_13416_));
 NAND3_X2 _22794_ (.A1(_13329_),
    .A2(_13286_),
    .A3(_13287_),
    .ZN(_13417_));
 NAND2_X1 _22795_ (.A1(_13399_),
    .A2(_13417_),
    .ZN(_13418_));
 MUX2_X1 _22796_ (.A(_13416_),
    .B(_13418_),
    .S(_13217_),
    .Z(_13419_));
 AOI221_X2 _22797_ (.A(_13404_),
    .B1(_13407_),
    .B2(_13410_),
    .C1(_13419_),
    .C2(_13324_),
    .ZN(_13420_));
 AOI222_X2 _22798_ (.A1(_13361_),
    .A2(_13322_),
    .B1(_13376_),
    .B2(_13392_),
    .C1(_13403_),
    .C2(_13420_),
    .ZN(_00080_));
 NAND2_X2 _22799_ (.A1(_13234_),
    .A2(_13274_),
    .ZN(_13421_));
 CLKBUF_X3 _22800_ (.A(_13298_),
    .Z(_13422_));
 AOI21_X1 _22801_ (.A(_13237_),
    .B1(_13283_),
    .B2(_13313_),
    .ZN(_13423_));
 MUX2_X1 _22802_ (.A(_13385_),
    .B(net176),
    .S(_13256_),
    .Z(_13424_));
 AOI21_X1 _22803_ (.A(_13423_),
    .B1(_13424_),
    .B2(_13238_),
    .ZN(_13425_));
 OAI21_X4 _22804_ (.A(_13332_),
    .B1(_13262_),
    .B2(_13263_),
    .ZN(_13426_));
 AOI21_X1 _22805_ (.A(_13218_),
    .B1(_13340_),
    .B2(_13426_),
    .ZN(_13427_));
 OAI21_X1 _22806_ (.A(_13298_),
    .B1(_13283_),
    .B2(_13223_),
    .ZN(_13428_));
 OAI22_X1 _22807_ (.A1(_13422_),
    .A2(_13425_),
    .B1(_13427_),
    .B2(_13428_),
    .ZN(_13429_));
 INV_X1 _22808_ (.A(_15012_),
    .ZN(_13430_));
 AOI21_X1 _22809_ (.A(_13347_),
    .B1(_13298_),
    .B2(_13430_),
    .ZN(_13431_));
 MUX2_X1 _22810_ (.A(_13289_),
    .B(_13415_),
    .S(_13223_),
    .Z(_13432_));
 AOI21_X1 _22811_ (.A(_13431_),
    .B1(_13432_),
    .B2(_13347_),
    .ZN(_13433_));
 OAI221_X1 _22812_ (.A(_13228_),
    .B1(_13421_),
    .B2(_13429_),
    .C1(_13433_),
    .C2(_13344_),
    .ZN(_13434_));
 AOI21_X1 _22813_ (.A(_13309_),
    .B1(_13283_),
    .B2(_13426_),
    .ZN(_13435_));
 INV_X1 _22814_ (.A(_13240_),
    .ZN(_13436_));
 NOR2_X1 _22815_ (.A1(_13436_),
    .A2(_13334_),
    .ZN(_13437_));
 AOI21_X2 _22816_ (.A(_14988_),
    .B1(_13286_),
    .B2(_13287_),
    .ZN(_13438_));
 NOR3_X1 _22817_ (.A1(_15011_),
    .A2(_13437_),
    .A3(_13438_),
    .ZN(_13439_));
 OAI21_X1 _22818_ (.A(_13379_),
    .B1(_13435_),
    .B2(_13439_),
    .ZN(_13440_));
 AND2_X1 _22819_ (.A1(_13255_),
    .A2(_13415_),
    .ZN(_13441_));
 OAI21_X1 _22820_ (.A(_13218_),
    .B1(_13334_),
    .B2(_13240_),
    .ZN(_13442_));
 AOI21_X2 _22821_ (.A(_13332_),
    .B1(_13286_),
    .B2(_13287_),
    .ZN(_13443_));
 NOR3_X4 _22822_ (.A1(_15002_),
    .A2(_13262_),
    .A3(_13263_),
    .ZN(_13444_));
 OR2_X1 _22823_ (.A1(_13443_),
    .A2(_13444_),
    .ZN(_13445_));
 OAI221_X1 _22824_ (.A(_13422_),
    .B1(_13441_),
    .B2(_13442_),
    .C1(_13445_),
    .C2(_15011_),
    .ZN(_13446_));
 AOI21_X1 _22825_ (.A(_13408_),
    .B1(_13440_),
    .B2(_13446_),
    .ZN(_13447_));
 NOR2_X4 _22826_ (.A1(net488),
    .A2(_13282_),
    .ZN(_13448_));
 NAND2_X2 _22827_ (.A1(_13197_),
    .A2(_13215_),
    .ZN(_13449_));
 AND2_X1 _22828_ (.A1(_13396_),
    .A2(_13449_),
    .ZN(_13450_));
 OAI21_X1 _22829_ (.A(_13396_),
    .B1(_13222_),
    .B2(_13385_),
    .ZN(_13451_));
 AOI221_X1 _22830_ (.A(_13297_),
    .B1(_13448_),
    .B2(_13450_),
    .C1(_13451_),
    .C2(_13346_),
    .ZN(_13452_));
 XNOR2_X1 _22831_ (.A(net1),
    .B(_13282_),
    .ZN(_13453_));
 AOI21_X1 _22832_ (.A(_13423_),
    .B1(_13453_),
    .B2(_13218_),
    .ZN(_13454_));
 NOR2_X1 _22833_ (.A1(_13378_),
    .A2(_13454_),
    .ZN(_13455_));
 NOR4_X2 _22834_ (.A1(_13364_),
    .A2(_13345_),
    .A3(_13452_),
    .A4(_13455_),
    .ZN(_13456_));
 NAND2_X1 _22835_ (.A1(_13301_),
    .A2(_13379_),
    .ZN(_13457_));
 NOR3_X1 _22836_ (.A1(_13348_),
    .A2(_13275_),
    .A3(_13339_),
    .ZN(_13458_));
 AOI21_X1 _22837_ (.A(_13302_),
    .B1(_13313_),
    .B2(_13458_),
    .ZN(_13459_));
 AOI21_X1 _22838_ (.A(_14995_),
    .B1(_13382_),
    .B2(_13383_),
    .ZN(_13460_));
 OAI22_X1 _22839_ (.A1(_13332_),
    .A2(_13288_),
    .B1(_13399_),
    .B2(_13178_),
    .ZN(_13461_));
 OAI21_X1 _22840_ (.A(_13276_),
    .B1(_13460_),
    .B2(_13461_),
    .ZN(_13462_));
 BUF_X4 _22841_ (.A(_13362_),
    .Z(_13463_));
 OAI21_X2 _22842_ (.A(_13305_),
    .B1(_13315_),
    .B2(_13316_),
    .ZN(_13464_));
 NAND3_X2 _22843_ (.A1(_14988_),
    .A2(_13286_),
    .A3(_13287_),
    .ZN(_13465_));
 AOI21_X1 _22844_ (.A(_13218_),
    .B1(_13464_),
    .B2(_13465_),
    .ZN(_13466_));
 NAND2_X1 _22845_ (.A1(_13463_),
    .A2(_13466_),
    .ZN(_13467_));
 NAND3_X1 _22846_ (.A1(_13459_),
    .A2(_13462_),
    .A3(_13467_),
    .ZN(_13468_));
 NAND2_X1 _22847_ (.A1(_13353_),
    .A2(_13237_),
    .ZN(_13469_));
 NAND2_X1 _22848_ (.A1(net175),
    .A2(_13222_),
    .ZN(_13470_));
 AOI21_X1 _22849_ (.A(_13346_),
    .B1(_13469_),
    .B2(_13470_),
    .ZN(_13471_));
 AOI21_X1 _22850_ (.A(_13409_),
    .B1(_13384_),
    .B2(_13178_),
    .ZN(_13472_));
 OAI221_X1 _22851_ (.A(_13236_),
    .B1(_13398_),
    .B2(_13471_),
    .C1(_13472_),
    .C2(_13276_),
    .ZN(_13473_));
 AND3_X1 _22852_ (.A1(_13457_),
    .A2(_13468_),
    .A3(_13473_),
    .ZN(_13474_));
 BUF_X32 _22853_ (.A(_13284_),
    .Z(_14987_));
 OAI21_X1 _22854_ (.A(_14987_),
    .B1(_13278_),
    .B2(_13339_),
    .ZN(_13475_));
 AOI21_X1 _22855_ (.A(_13363_),
    .B1(_13449_),
    .B2(_13475_),
    .ZN(_13476_));
 NOR2_X1 _22856_ (.A1(_13364_),
    .A2(_13298_),
    .ZN(_13477_));
 AND2_X1 _22857_ (.A1(_13417_),
    .A2(_13464_),
    .ZN(_13478_));
 NAND2_X1 _22858_ (.A1(_13222_),
    .A2(_13362_),
    .ZN(_13479_));
 OAI21_X1 _22859_ (.A(_13477_),
    .B1(_13478_),
    .B2(_13479_),
    .ZN(_13480_));
 NOR3_X4 _22860_ (.A1(_13197_),
    .A2(_13315_),
    .A3(_13316_),
    .ZN(_13481_));
 OAI21_X1 _22861_ (.A(_13481_),
    .B1(_13463_),
    .B2(net178),
    .ZN(_13482_));
 AOI21_X1 _22862_ (.A(_13338_),
    .B1(_13399_),
    .B2(_13482_),
    .ZN(_13483_));
 NOR3_X1 _22863_ (.A1(_13476_),
    .A2(_13480_),
    .A3(_13483_),
    .ZN(_13484_));
 NOR2_X1 _22864_ (.A1(_13348_),
    .A2(_13416_),
    .ZN(_13485_));
 AND3_X1 _22865_ (.A1(_13222_),
    .A2(_13426_),
    .A3(_13417_),
    .ZN(_13486_));
 AOI21_X1 _22866_ (.A(_13337_),
    .B1(_13257_),
    .B2(net175),
    .ZN(_13487_));
 OAI21_X1 _22867_ (.A(_13362_),
    .B1(_13328_),
    .B2(net177),
    .ZN(_13488_));
 NAND2_X1 _22868_ (.A1(_13177_),
    .A2(_14995_),
    .ZN(_13489_));
 NOR2_X1 _22869_ (.A1(_13257_),
    .A2(_13489_),
    .ZN(_13490_));
 OAI33_X1 _22870_ (.A1(_13463_),
    .A2(_13485_),
    .A3(_13486_),
    .B1(_13487_),
    .B2(_13488_),
    .B3(_13490_),
    .ZN(_13491_));
 NOR3_X1 _22871_ (.A1(_13371_),
    .A2(_13422_),
    .A3(_13491_),
    .ZN(_13492_));
 OAI33_X1 _22872_ (.A1(_13434_),
    .A2(_13447_),
    .A3(_13456_),
    .B1(_13492_),
    .B2(_13484_),
    .B3(_13474_),
    .ZN(_00081_));
 NOR2_X2 _22873_ (.A1(_13274_),
    .A2(_13377_),
    .ZN(_13493_));
 AOI21_X1 _22874_ (.A(_13348_),
    .B1(_13426_),
    .B2(_13465_),
    .ZN(_13494_));
 BUF_X4 _22875_ (.A(_13282_),
    .Z(_13495_));
 AOI211_X2 _22876_ (.A(_13216_),
    .B(_13304_),
    .C1(_13495_),
    .C2(net176),
    .ZN(_13496_));
 NOR3_X1 _22877_ (.A1(_13371_),
    .A2(_13494_),
    .A3(_13496_),
    .ZN(_13497_));
 INV_X1 _22878_ (.A(_15016_),
    .ZN(_13498_));
 AOI221_X2 _22879_ (.A(_13234_),
    .B1(_13448_),
    .B2(_13449_),
    .C1(_13346_),
    .C2(_13498_),
    .ZN(_13499_));
 OAI21_X1 _22880_ (.A(_13493_),
    .B1(_13497_),
    .B2(_13499_),
    .ZN(_13500_));
 NAND2_X2 _22881_ (.A1(_13274_),
    .A2(_13297_),
    .ZN(_13501_));
 NAND2_X1 _22882_ (.A1(_13234_),
    .A2(_13381_),
    .ZN(_13502_));
 NAND3_X1 _22883_ (.A1(_13237_),
    .A2(_13323_),
    .A3(_13481_),
    .ZN(_13503_));
 AOI21_X1 _22884_ (.A(_13284_),
    .B1(_13502_),
    .B2(_13503_),
    .ZN(_13504_));
 AOI21_X1 _22885_ (.A(_13234_),
    .B1(_13256_),
    .B2(_15007_),
    .ZN(_13505_));
 AOI21_X4 _22886_ (.A(_13197_),
    .B1(_13249_),
    .B2(_13253_),
    .ZN(_13506_));
 AOI22_X1 _22887_ (.A1(_15012_),
    .A2(_13495_),
    .B1(_13506_),
    .B2(net133),
    .ZN(_13507_));
 AOI21_X1 _22888_ (.A(_13505_),
    .B1(_13507_),
    .B2(_13235_),
    .ZN(_13508_));
 OR3_X1 _22889_ (.A1(_13501_),
    .A2(_13504_),
    .A3(_13508_),
    .ZN(_13509_));
 AND3_X1 _22890_ (.A1(_13301_),
    .A2(_13500_),
    .A3(_13509_),
    .ZN(_13510_));
 NAND3_X1 _22891_ (.A1(_14992_),
    .A2(_13223_),
    .A3(_13399_),
    .ZN(_13511_));
 NAND2_X1 _22892_ (.A1(_14995_),
    .A2(_13222_),
    .ZN(_13512_));
 NAND3_X1 _22893_ (.A1(net141),
    .A2(_13334_),
    .A3(_13512_),
    .ZN(_13513_));
 NAND2_X1 _22894_ (.A1(_13511_),
    .A2(_13513_),
    .ZN(_13514_));
 MUX2_X1 _22895_ (.A(_13222_),
    .B(_13257_),
    .S(_13177_),
    .Z(_13515_));
 OAI21_X1 _22896_ (.A(_13235_),
    .B1(_13515_),
    .B2(net611),
    .ZN(_13516_));
 NOR2_X1 _22897_ (.A1(_14990_),
    .A2(_14993_),
    .ZN(_13517_));
 AOI221_X2 _22898_ (.A(_13215_),
    .B1(_13255_),
    .B2(_13517_),
    .C1(_13339_),
    .C2(_13176_),
    .ZN(_13518_));
 AOI21_X1 _22899_ (.A(_13348_),
    .B1(_13346_),
    .B2(_13289_),
    .ZN(_13519_));
 NAND2_X1 _22900_ (.A1(_13334_),
    .A2(_13415_),
    .ZN(_13520_));
 AOI21_X1 _22901_ (.A(_13518_),
    .B1(_13519_),
    .B2(_13520_),
    .ZN(_13521_));
 OAI221_X1 _22902_ (.A(_13363_),
    .B1(_13514_),
    .B2(_13516_),
    .C1(_13521_),
    .C2(_13364_),
    .ZN(_13522_));
 OAI221_X1 _22903_ (.A(_13393_),
    .B1(_13396_),
    .B2(_14987_),
    .C1(_13338_),
    .C2(_13353_),
    .ZN(_13523_));
 AOI21_X1 _22904_ (.A(_13421_),
    .B1(_13347_),
    .B2(_15009_),
    .ZN(_13524_));
 NAND3_X1 _22905_ (.A1(_13338_),
    .A2(_13426_),
    .A3(_13465_),
    .ZN(_13525_));
 AOI21_X1 _22906_ (.A(_13344_),
    .B1(_13278_),
    .B2(net540),
    .ZN(_13526_));
 AOI22_X1 _22907_ (.A1(_13523_),
    .A2(_13524_),
    .B1(_13525_),
    .B2(_13526_),
    .ZN(_13527_));
 NAND3_X1 _22908_ (.A1(_13379_),
    .A2(_13522_),
    .A3(_13527_),
    .ZN(_13528_));
 NOR2_X1 _22909_ (.A1(_13234_),
    .A2(_13362_),
    .ZN(_13529_));
 AOI21_X4 _22910_ (.A(_14998_),
    .B1(_13249_),
    .B2(_13253_),
    .ZN(_13530_));
 NOR3_X1 _22911_ (.A1(_13218_),
    .A2(_13481_),
    .A3(_13530_),
    .ZN(_13531_));
 NOR3_X1 _22912_ (.A1(_13337_),
    .A2(_13448_),
    .A3(_13444_),
    .ZN(_13532_));
 NOR3_X1 _22913_ (.A1(_13408_),
    .A2(_13531_),
    .A3(_13532_),
    .ZN(_13533_));
 NOR3_X1 _22914_ (.A1(_13337_),
    .A2(_13406_),
    .A3(_13443_),
    .ZN(_13534_));
 NOR3_X1 _22915_ (.A1(_13405_),
    .A2(_13481_),
    .A3(_13237_),
    .ZN(_13535_));
 AOI21_X2 _22916_ (.A(_13217_),
    .B1(_13399_),
    .B2(_13372_),
    .ZN(_13536_));
 AOI21_X1 _22917_ (.A(_13240_),
    .B1(_13286_),
    .B2(_13287_),
    .ZN(_13537_));
 NOR3_X1 _22918_ (.A1(_13222_),
    .A2(_13537_),
    .A3(_13366_),
    .ZN(_13538_));
 OAI33_X1 _22919_ (.A1(_13463_),
    .A2(_13534_),
    .A3(_13535_),
    .B1(_13536_),
    .B2(_13538_),
    .B3(_13235_),
    .ZN(_13539_));
 OR3_X1 _22920_ (.A1(_13539_),
    .A2(_13533_),
    .A3(_13529_),
    .ZN(_13540_));
 NAND2_X1 _22921_ (.A1(_13228_),
    .A2(_13379_),
    .ZN(_13541_));
 NOR4_X1 _22922_ (.A1(_14987_),
    .A2(_13348_),
    .A3(_13506_),
    .A4(_13339_),
    .ZN(_13542_));
 NOR2_X1 _22923_ (.A1(net175),
    .A2(_13328_),
    .ZN(_13543_));
 NOR3_X1 _22924_ (.A1(_13344_),
    .A2(_13542_),
    .A3(_13543_),
    .ZN(_13544_));
 NOR2_X1 _22925_ (.A1(_13541_),
    .A2(_13544_),
    .ZN(_13545_));
 NOR2_X4 _22926_ (.A1(net495),
    .A2(_13220_),
    .ZN(_13546_));
 AND2_X1 _22927_ (.A1(_13277_),
    .A2(_13282_),
    .ZN(_13547_));
 NOR3_X1 _22928_ (.A1(_13217_),
    .A2(_13448_),
    .A3(_13547_),
    .ZN(_13548_));
 NOR3_X1 _22929_ (.A1(_13421_),
    .A2(_13546_),
    .A3(_13548_),
    .ZN(_13549_));
 NOR3_X1 _22930_ (.A1(_13217_),
    .A2(_13265_),
    .A3(_13368_),
    .ZN(_13550_));
 AOI21_X2 _22931_ (.A(_13329_),
    .B1(_13286_),
    .B2(_13287_),
    .ZN(_13551_));
 NOR3_X1 _22932_ (.A1(_13309_),
    .A2(_13551_),
    .A3(_13306_),
    .ZN(_13552_));
 OR2_X1 _22933_ (.A1(_13550_),
    .A2(_13552_),
    .ZN(_13553_));
 NOR3_X1 _22934_ (.A1(_13216_),
    .A2(_13506_),
    .A3(_13406_),
    .ZN(_13554_));
 NOR3_X2 _22935_ (.A1(_13309_),
    .A2(_13551_),
    .A3(_13444_),
    .ZN(_13555_));
 NOR3_X1 _22936_ (.A1(_13323_),
    .A2(_13554_),
    .A3(_13555_),
    .ZN(_13556_));
 NOR3_X4 _22937_ (.A1(_13214_),
    .A2(_13262_),
    .A3(_13263_),
    .ZN(_13557_));
 OAI21_X1 _22938_ (.A(_13399_),
    .B1(_13255_),
    .B2(_13356_),
    .ZN(_13558_));
 AOI221_X2 _22939_ (.A(_13325_),
    .B1(_13557_),
    .B2(net540),
    .C1(_13558_),
    .C2(_13216_),
    .ZN(_13559_));
 AOI21_X1 _22940_ (.A(_13556_),
    .B1(_13559_),
    .B2(_13323_),
    .ZN(_13560_));
 AOI221_X2 _22941_ (.A(_13549_),
    .B1(_13553_),
    .B2(_13529_),
    .C1(_13560_),
    .C2(_13463_),
    .ZN(_13561_));
 NOR2_X1 _22942_ (.A1(_13301_),
    .A2(_13379_),
    .ZN(_13562_));
 AOI222_X2 _22943_ (.A1(_13510_),
    .A2(_13528_),
    .B1(_13545_),
    .B2(_13540_),
    .C1(_13561_),
    .C2(_13562_),
    .ZN(_00082_));
 NAND2_X1 _22944_ (.A1(_13236_),
    .A2(_13378_),
    .ZN(_13563_));
 NOR2_X1 _22945_ (.A1(_13289_),
    .A2(_13393_),
    .ZN(_13564_));
 NOR3_X1 _22946_ (.A1(_15011_),
    .A2(_13564_),
    .A3(_13438_),
    .ZN(_13565_));
 NOR3_X1 _22947_ (.A1(_13338_),
    .A2(_13339_),
    .A3(_13405_),
    .ZN(_13566_));
 OAI21_X1 _22948_ (.A(_13363_),
    .B1(_13565_),
    .B2(_13566_),
    .ZN(_13567_));
 NAND2_X1 _22949_ (.A1(_13356_),
    .A2(_13393_),
    .ZN(_13568_));
 NAND3_X1 _22950_ (.A1(_15004_),
    .A2(_13372_),
    .A3(_13568_),
    .ZN(_13569_));
 OR3_X1 _22951_ (.A1(_13338_),
    .A2(_13551_),
    .A3(_13368_),
    .ZN(_13570_));
 NAND3_X1 _22952_ (.A1(_13345_),
    .A2(_13569_),
    .A3(_13570_),
    .ZN(_13571_));
 AOI21_X1 _22953_ (.A(_13563_),
    .B1(_13567_),
    .B2(_13571_),
    .ZN(_13572_));
 INV_X1 _22954_ (.A(_13289_),
    .ZN(_13573_));
 OAI221_X1 _22955_ (.A(_13275_),
    .B1(_13288_),
    .B2(_13353_),
    .C1(_13328_),
    .C2(_13573_),
    .ZN(_13574_));
 OAI22_X1 _22956_ (.A1(_14995_),
    .A2(_13382_),
    .B1(_13512_),
    .B2(_13393_),
    .ZN(_13575_));
 AOI21_X1 _22957_ (.A(_13574_),
    .B1(_13575_),
    .B2(net178),
    .ZN(_13576_));
 OAI221_X1 _22958_ (.A(_13463_),
    .B1(_13264_),
    .B2(_13178_),
    .C1(_13288_),
    .C2(_13573_),
    .ZN(_13577_));
 OAI21_X1 _22959_ (.A(_13379_),
    .B1(_13536_),
    .B2(_13577_),
    .ZN(_13578_));
 NOR3_X1 _22960_ (.A1(_13302_),
    .A2(_13576_),
    .A3(_13578_),
    .ZN(_13579_));
 NOR3_X2 _22961_ (.A1(_13228_),
    .A2(_13235_),
    .A3(_13378_),
    .ZN(_13580_));
 NOR4_X1 _22962_ (.A1(net133),
    .A2(_13221_),
    .A3(_13299_),
    .A4(_13282_),
    .ZN(_13581_));
 NAND2_X1 _22963_ (.A1(_13217_),
    .A2(_13274_),
    .ZN(_13582_));
 AOI221_X1 _22964_ (.A(_13581_),
    .B1(_13582_),
    .B2(_13443_),
    .C1(_13362_),
    .C2(_13381_),
    .ZN(_13583_));
 NOR3_X1 _22965_ (.A1(_13219_),
    .A2(_13217_),
    .A3(_13274_),
    .ZN(_13584_));
 NAND2_X1 _22966_ (.A1(_13219_),
    .A2(_13274_),
    .ZN(_13585_));
 NOR2_X1 _22967_ (.A1(net133),
    .A2(_13288_),
    .ZN(_13586_));
 NOR2_X2 _22968_ (.A1(_13219_),
    .A2(_13215_),
    .ZN(_13587_));
 NOR2_X1 _22969_ (.A1(_13300_),
    .A2(_13587_),
    .ZN(_13588_));
 AOI221_X2 _22970_ (.A(_13584_),
    .B1(_13585_),
    .B2(_13586_),
    .C1(_13588_),
    .C2(_13368_),
    .ZN(_13589_));
 NAND3_X1 _22971_ (.A1(_13580_),
    .A2(_13583_),
    .A3(_13589_),
    .ZN(_13590_));
 OAI21_X1 _22972_ (.A(_13273_),
    .B1(_13197_),
    .B2(net173),
    .ZN(_13591_));
 NOR2_X1 _22973_ (.A1(net612),
    .A2(_13383_),
    .ZN(_13592_));
 OAI21_X1 _22974_ (.A(_13449_),
    .B1(_13339_),
    .B2(net176),
    .ZN(_13593_));
 AOI221_X1 _22975_ (.A(_13378_),
    .B1(_13591_),
    .B2(_13592_),
    .C1(_13593_),
    .C2(_13274_),
    .ZN(_13594_));
 AOI21_X1 _22976_ (.A(_13547_),
    .B1(_13393_),
    .B2(net175),
    .ZN(_13595_));
 NAND2_X1 _22977_ (.A1(_13216_),
    .A2(_13299_),
    .ZN(_13596_));
 OAI221_X1 _22978_ (.A(_13594_),
    .B1(_13595_),
    .B2(_13596_),
    .C1(_14987_),
    .C2(_13328_),
    .ZN(_13597_));
 OAI21_X1 _22979_ (.A(_13590_),
    .B1(_13597_),
    .B2(_13302_),
    .ZN(_13598_));
 NOR2_X2 _22980_ (.A1(_13196_),
    .A2(_13383_),
    .ZN(_13599_));
 AND2_X1 _22981_ (.A1(_13277_),
    .A2(_13377_),
    .ZN(_13600_));
 NOR2_X2 _22982_ (.A1(_13278_),
    .A2(_13557_),
    .ZN(_13601_));
 AOI221_X2 _22983_ (.A(_13299_),
    .B1(_13377_),
    .B2(_13599_),
    .C1(_13600_),
    .C2(_13601_),
    .ZN(_13602_));
 OR2_X4 _22984_ (.A1(_14993_),
    .A2(_14990_),
    .ZN(_13603_));
 OAI21_X4 _22985_ (.A(_13603_),
    .B1(_13263_),
    .B2(_13262_),
    .ZN(_13604_));
 AND2_X2 _22986_ (.A1(_13604_),
    .A2(_13372_),
    .ZN(_13605_));
 OAI21_X1 _22987_ (.A(_13283_),
    .B1(_13281_),
    .B2(_13355_),
    .ZN(_13606_));
 MUX2_X1 _22988_ (.A(_13605_),
    .B(_13606_),
    .S(_13215_),
    .Z(_13607_));
 OAI22_X1 _22989_ (.A1(_13436_),
    .A2(_13281_),
    .B1(_13333_),
    .B2(_13296_),
    .ZN(_13608_));
 AOI21_X2 _22990_ (.A(_13273_),
    .B1(_13608_),
    .B2(_13221_),
    .ZN(_13609_));
 OAI21_X1 _22991_ (.A(_13426_),
    .B1(_13254_),
    .B2(_14996_),
    .ZN(_13610_));
 AOI22_X2 _22992_ (.A1(net174),
    .A2(_13557_),
    .B1(_13610_),
    .B2(_13215_),
    .ZN(_13611_));
 AOI221_X2 _22993_ (.A(_13234_),
    .B1(_13607_),
    .B2(_13602_),
    .C1(_13609_),
    .C2(_13611_),
    .ZN(_13612_));
 OAI21_X1 _22994_ (.A(_13378_),
    .B1(_13602_),
    .B2(_13609_),
    .ZN(_13613_));
 NOR2_X4 _22995_ (.A1(_13273_),
    .A2(_13297_),
    .ZN(_13614_));
 OAI21_X1 _22996_ (.A(_13220_),
    .B1(_13306_),
    .B2(_13530_),
    .ZN(_13615_));
 OAI21_X1 _22997_ (.A(_13264_),
    .B1(_13255_),
    .B2(_13356_),
    .ZN(_13616_));
 OAI21_X1 _22998_ (.A(_13615_),
    .B1(_13616_),
    .B2(_13221_),
    .ZN(_13617_));
 NOR2_X1 _22999_ (.A1(_13256_),
    .A2(_13357_),
    .ZN(_13618_));
 NAND2_X1 _23000_ (.A1(_13299_),
    .A2(_13297_),
    .ZN(_13619_));
 NOR2_X1 _23001_ (.A1(_13619_),
    .A2(_13587_),
    .ZN(_13620_));
 AOI221_X2 _23002_ (.A(_13323_),
    .B1(_13614_),
    .B2(_13617_),
    .C1(_13618_),
    .C2(_13620_),
    .ZN(_13621_));
 OAI21_X1 _23003_ (.A(_13216_),
    .B1(_13256_),
    .B2(_13573_),
    .ZN(_13622_));
 OR2_X1 _23004_ (.A1(_13622_),
    .A2(_13530_),
    .ZN(_13623_));
 NOR2_X1 _23005_ (.A1(_13501_),
    .A2(_13518_),
    .ZN(_13624_));
 OAI21_X1 _23006_ (.A(_14995_),
    .B1(_13237_),
    .B2(_13368_),
    .ZN(_13625_));
 NAND2_X1 _23007_ (.A1(_13273_),
    .A2(_13377_),
    .ZN(_13626_));
 AOI221_X2 _23008_ (.A(_13626_),
    .B1(_13317_),
    .B2(net173),
    .C1(_13385_),
    .C2(_13381_),
    .ZN(_13627_));
 AOI22_X2 _23009_ (.A1(_13623_),
    .A2(_13624_),
    .B1(_13625_),
    .B2(_13627_),
    .ZN(_13628_));
 AOI221_X2 _23010_ (.A(_13301_),
    .B1(_13612_),
    .B2(_13613_),
    .C1(_13621_),
    .C2(_13628_),
    .ZN(_13629_));
 NOR4_X2 _23011_ (.A1(_13579_),
    .A2(_13629_),
    .A3(_13598_),
    .A4(_13572_),
    .ZN(_00083_));
 NAND2_X1 _23012_ (.A1(_15000_),
    .A2(_13346_),
    .ZN(_13630_));
 OAI21_X1 _23013_ (.A(_13630_),
    .B1(_13469_),
    .B2(_13347_),
    .ZN(_13631_));
 AOI21_X1 _23014_ (.A(_15004_),
    .B1(_13399_),
    .B2(_13465_),
    .ZN(_13632_));
 OAI221_X2 _23015_ (.A(_13422_),
    .B1(_13383_),
    .B2(_13240_),
    .C1(_14987_),
    .C2(_13264_),
    .ZN(_13633_));
 OAI221_X2 _23016_ (.A(_13345_),
    .B1(_13422_),
    .B2(_13631_),
    .C1(_13632_),
    .C2(_13633_),
    .ZN(_13634_));
 AND2_X1 _23017_ (.A1(_13347_),
    .A2(_13350_),
    .ZN(_13635_));
 OAI21_X1 _23018_ (.A(_15004_),
    .B1(_13635_),
    .B2(_13448_),
    .ZN(_13636_));
 NAND3_X1 _23019_ (.A1(_13279_),
    .A2(_13614_),
    .A3(_13636_),
    .ZN(_13637_));
 NAND2_X1 _23020_ (.A1(_13228_),
    .A2(_13371_),
    .ZN(_13638_));
 AND3_X1 _23021_ (.A1(_13279_),
    .A2(_13340_),
    .A3(_13493_),
    .ZN(_13639_));
 OAI21_X1 _23022_ (.A(_15004_),
    .B1(_13506_),
    .B2(_13368_),
    .ZN(_13640_));
 AOI21_X1 _23023_ (.A(_13638_),
    .B1(_13639_),
    .B2(_13640_),
    .ZN(_13641_));
 NAND3_X1 _23024_ (.A1(_13634_),
    .A2(_13637_),
    .A3(_13641_),
    .ZN(_13642_));
 AOI21_X1 _23025_ (.A(_13197_),
    .B1(_13216_),
    .B2(_13273_),
    .ZN(_13643_));
 OAI221_X2 _23026_ (.A(_13495_),
    .B1(_13643_),
    .B2(net133),
    .C1(_13219_),
    .C2(_13217_),
    .ZN(_13644_));
 NAND2_X1 _23027_ (.A1(net176),
    .A2(_13309_),
    .ZN(_13645_));
 OAI221_X2 _23028_ (.A(_13256_),
    .B1(_13596_),
    .B2(_13385_),
    .C1(_13645_),
    .C2(_13300_),
    .ZN(_13646_));
 NAND2_X1 _23029_ (.A1(_13274_),
    .A2(_13506_),
    .ZN(_13647_));
 NAND2_X1 _23030_ (.A1(_13479_),
    .A2(_13647_),
    .ZN(_13648_));
 AOI221_X1 _23031_ (.A(_13404_),
    .B1(_13644_),
    .B2(_13646_),
    .C1(_13648_),
    .C2(net141),
    .ZN(_13649_));
 NOR2_X1 _23032_ (.A1(_13228_),
    .A2(_13298_),
    .ZN(_13650_));
 OAI21_X2 _23033_ (.A(_13277_),
    .B1(_13315_),
    .B2(_13316_),
    .ZN(_13651_));
 AND2_X1 _23034_ (.A1(_13237_),
    .A2(_13651_),
    .ZN(_13652_));
 OAI21_X1 _23035_ (.A(_13463_),
    .B1(_13258_),
    .B2(_13652_),
    .ZN(_13653_));
 OAI21_X2 _23036_ (.A(_13237_),
    .B1(_13495_),
    .B2(_13284_),
    .ZN(_13654_));
 NOR2_X1 _23037_ (.A1(_13385_),
    .A2(_13257_),
    .ZN(_13655_));
 OAI21_X1 _23038_ (.A(_13588_),
    .B1(_13654_),
    .B2(_13655_),
    .ZN(_13656_));
 AND3_X1 _23039_ (.A1(_13650_),
    .A2(_13653_),
    .A3(_13656_),
    .ZN(_13657_));
 NOR3_X1 _23040_ (.A1(_13236_),
    .A2(_13649_),
    .A3(_13657_),
    .ZN(_13658_));
 NAND2_X1 _23041_ (.A1(_13300_),
    .A2(_13377_),
    .ZN(_13659_));
 AOI21_X1 _23042_ (.A(_13309_),
    .B1(_13417_),
    .B2(_13464_),
    .ZN(_13660_));
 AOI21_X1 _23043_ (.A(_13660_),
    .B1(_13337_),
    .B2(_13277_),
    .ZN(_13661_));
 OAI21_X1 _23044_ (.A(_13371_),
    .B1(_13659_),
    .B2(_13661_),
    .ZN(_13662_));
 NOR2_X1 _23045_ (.A1(_13306_),
    .A2(_13530_),
    .ZN(_13663_));
 NOR2_X1 _23046_ (.A1(_13215_),
    .A2(_13444_),
    .ZN(_13664_));
 NAND2_X2 _23047_ (.A1(net173),
    .A2(_13506_),
    .ZN(_13665_));
 AOI221_X1 _23048_ (.A(_13297_),
    .B1(_13663_),
    .B2(_13215_),
    .C1(_13664_),
    .C2(_13665_),
    .ZN(_13666_));
 NOR2_X1 _23049_ (.A1(_13197_),
    .A2(_13214_),
    .ZN(_13667_));
 NAND2_X1 _23050_ (.A1(net173),
    .A2(_13667_),
    .ZN(_13668_));
 NOR2_X1 _23051_ (.A1(_13255_),
    .A2(_13546_),
    .ZN(_13669_));
 NAND2_X1 _23052_ (.A1(_13385_),
    .A2(_13220_),
    .ZN(_13670_));
 OAI21_X1 _23053_ (.A(_13670_),
    .B1(_13220_),
    .B2(_13175_),
    .ZN(_13671_));
 AOI221_X2 _23054_ (.A(_13299_),
    .B1(_13668_),
    .B2(_13669_),
    .C1(_13671_),
    .C2(_13255_),
    .ZN(_13672_));
 AOI21_X2 _23055_ (.A(_13666_),
    .B1(_13672_),
    .B2(_13297_),
    .ZN(_13673_));
 AOI21_X2 _23056_ (.A(_13444_),
    .B1(_13256_),
    .B2(net1),
    .ZN(_13674_));
 NOR3_X2 _23057_ (.A1(_13329_),
    .A2(_13315_),
    .A3(_13316_),
    .ZN(_13675_));
 NOR2_X1 _23058_ (.A1(_13217_),
    .A2(_13675_),
    .ZN(_13676_));
 AOI22_X1 _23059_ (.A1(_13218_),
    .A2(_13674_),
    .B1(_13676_),
    .B2(_13665_),
    .ZN(_13677_));
 NOR2_X1 _23060_ (.A1(_13672_),
    .A2(_13677_),
    .ZN(_13678_));
 AOI221_X2 _23061_ (.A(_13662_),
    .B1(_13673_),
    .B2(_13276_),
    .C1(_13298_),
    .C2(_13678_),
    .ZN(_13679_));
 NOR2_X1 _23062_ (.A1(_13301_),
    .A2(_13371_),
    .ZN(_13680_));
 INV_X1 _23063_ (.A(_13680_),
    .ZN(_13681_));
 NOR2_X1 _23064_ (.A1(_15004_),
    .A2(_13276_),
    .ZN(_13682_));
 AOI21_X1 _23065_ (.A(_13422_),
    .B1(_13441_),
    .B2(_13682_),
    .ZN(_13683_));
 AOI21_X1 _23066_ (.A(_13675_),
    .B1(_13415_),
    .B2(_13393_),
    .ZN(_13684_));
 OAI21_X1 _23067_ (.A(_15004_),
    .B1(_13363_),
    .B2(_13684_),
    .ZN(_13685_));
 MUX2_X1 _23068_ (.A(net611),
    .B(_13240_),
    .S(_13362_),
    .Z(_13686_));
 OAI21_X1 _23069_ (.A(_13647_),
    .B1(_13686_),
    .B2(_13393_),
    .ZN(_13687_));
 OAI21_X1 _23070_ (.A(_13685_),
    .B1(_13687_),
    .B2(_15004_),
    .ZN(_13688_));
 OAI21_X1 _23071_ (.A(_13313_),
    .B1(_13257_),
    .B2(_14988_),
    .ZN(_13689_));
 MUX2_X1 _23072_ (.A(_13453_),
    .B(_13689_),
    .S(_13337_),
    .Z(_13690_));
 AOI22_X1 _23073_ (.A1(_13223_),
    .A2(_13283_),
    .B1(_13317_),
    .B2(_13356_),
    .ZN(_13691_));
 MUX2_X1 _23074_ (.A(_13690_),
    .B(_13691_),
    .S(_13276_),
    .Z(_13692_));
 AOI22_X1 _23075_ (.A1(_13683_),
    .A2(_13688_),
    .B1(_13692_),
    .B2(_13422_),
    .ZN(_13693_));
 OAI221_X1 _23076_ (.A(_13642_),
    .B1(_13658_),
    .B2(_13679_),
    .C1(_13681_),
    .C2(_13693_),
    .ZN(_00084_));
 OAI21_X1 _23077_ (.A(_13377_),
    .B1(_13327_),
    .B2(_13603_),
    .ZN(_13694_));
 NAND2_X1 _23078_ (.A1(_13356_),
    .A2(_13216_),
    .ZN(_13695_));
 AOI22_X2 _23079_ (.A1(net540),
    .A2(_13317_),
    .B1(_13695_),
    .B2(_13256_),
    .ZN(_13696_));
 AOI221_X1 _23080_ (.A(_13694_),
    .B1(_13696_),
    .B2(_13300_),
    .C1(_13366_),
    .C2(_13450_),
    .ZN(_13697_));
 AOI221_X2 _23081_ (.A(_13501_),
    .B1(_13557_),
    .B2(_13415_),
    .C1(_13289_),
    .C2(_13257_),
    .ZN(_13698_));
 NOR2_X1 _23082_ (.A1(_13697_),
    .A2(_13698_),
    .ZN(_13699_));
 AOI21_X1 _23083_ (.A(_13276_),
    .B1(_13378_),
    .B2(_13696_),
    .ZN(_13700_));
 OAI21_X1 _23084_ (.A(_13223_),
    .B1(_13306_),
    .B2(_13443_),
    .ZN(_13701_));
 AOI21_X1 _23085_ (.A(_13304_),
    .B1(_13282_),
    .B2(_13355_),
    .ZN(_13702_));
 OAI21_X1 _23086_ (.A(_13701_),
    .B1(_13702_),
    .B2(_13338_),
    .ZN(_13703_));
 OAI21_X1 _23087_ (.A(_13700_),
    .B1(_13703_),
    .B2(_13379_),
    .ZN(_13704_));
 AOI21_X1 _23088_ (.A(_13638_),
    .B1(_13699_),
    .B2(_13704_),
    .ZN(_13705_));
 MUX2_X1 _23089_ (.A(_13356_),
    .B(_13176_),
    .S(_13281_),
    .Z(_13706_));
 AOI21_X1 _23090_ (.A(_13314_),
    .B1(_13216_),
    .B2(_13706_),
    .ZN(_13707_));
 AOI21_X1 _23091_ (.A(_13377_),
    .B1(_13278_),
    .B2(_13197_),
    .ZN(_13708_));
 AOI221_X2 _23092_ (.A(_13362_),
    .B1(_13707_),
    .B2(_13377_),
    .C1(_13708_),
    .C2(_13615_),
    .ZN(_13709_));
 NAND2_X1 _23093_ (.A1(_13223_),
    .A2(_13417_),
    .ZN(_13710_));
 AOI21_X1 _23094_ (.A(_13619_),
    .B1(_13710_),
    .B2(_13665_),
    .ZN(_13711_));
 NAND2_X1 _23095_ (.A1(_13277_),
    .A2(_13317_),
    .ZN(_13712_));
 AND4_X1 _23096_ (.A1(_13285_),
    .A2(_13313_),
    .A3(_13614_),
    .A4(_13712_),
    .ZN(_13713_));
 NOR4_X1 _23097_ (.A1(_13302_),
    .A2(_13709_),
    .A3(_13711_),
    .A4(_13713_),
    .ZN(_13714_));
 AOI21_X1 _23098_ (.A(_13348_),
    .B1(_13311_),
    .B2(_13464_),
    .ZN(_13715_));
 OAI21_X1 _23099_ (.A(_13362_),
    .B1(_13383_),
    .B2(net177),
    .ZN(_13716_));
 AOI21_X1 _23100_ (.A(_13438_),
    .B1(_13495_),
    .B2(_13355_),
    .ZN(_13717_));
 OAI22_X1 _23101_ (.A1(_13353_),
    .A2(_13328_),
    .B1(_13717_),
    .B2(_13348_),
    .ZN(_13718_));
 OAI221_X1 _23102_ (.A(_13580_),
    .B1(_13715_),
    .B2(_13716_),
    .C1(_13718_),
    .C2(_13463_),
    .ZN(_13719_));
 NOR2_X2 _23103_ (.A1(_13300_),
    .A2(_13495_),
    .ZN(_13720_));
 OAI21_X1 _23104_ (.A(_13284_),
    .B1(_13557_),
    .B2(_13720_),
    .ZN(_13721_));
 AOI22_X1 _23105_ (.A1(_13289_),
    .A2(_13278_),
    .B1(_13557_),
    .B2(_14986_),
    .ZN(_13722_));
 NAND2_X1 _23106_ (.A1(_13300_),
    .A2(_13495_),
    .ZN(_13723_));
 MUX2_X1 _23107_ (.A(_13256_),
    .B(_13327_),
    .S(_13299_),
    .Z(_13724_));
 MUX2_X1 _23108_ (.A(_13723_),
    .B(_13724_),
    .S(_13177_),
    .Z(_13725_));
 OAI221_X1 _23109_ (.A(_13721_),
    .B1(_13722_),
    .B2(_13276_),
    .C1(_14986_),
    .C2(_13725_),
    .ZN(_13726_));
 OAI21_X1 _23110_ (.A(_13719_),
    .B1(_13726_),
    .B2(_13563_),
    .ZN(_13727_));
 AOI221_X2 _23111_ (.A(_13409_),
    .B1(_13441_),
    .B2(_13221_),
    .C1(_13384_),
    .C2(_13219_),
    .ZN(_13728_));
 NOR2_X1 _23112_ (.A1(_13501_),
    .A2(_13728_),
    .ZN(_13729_));
 NOR2_X1 _23113_ (.A1(_13221_),
    .A2(_13406_),
    .ZN(_13730_));
 NOR2_X1 _23114_ (.A1(_13368_),
    .A2(_13405_),
    .ZN(_13731_));
 AOI221_X1 _23115_ (.A(_13659_),
    .B1(_13730_),
    .B2(_13665_),
    .C1(_13731_),
    .C2(_13309_),
    .ZN(_13732_));
 OAI221_X1 _23116_ (.A(_13493_),
    .B1(_13702_),
    .B2(_13222_),
    .C1(_13415_),
    .C2(_13383_),
    .ZN(_13733_));
 NAND2_X1 _23117_ (.A1(net176),
    .A2(_13495_),
    .ZN(_13734_));
 AOI21_X1 _23118_ (.A(_13599_),
    .B1(_13734_),
    .B2(_14986_),
    .ZN(_13735_));
 OAI21_X1 _23119_ (.A(_13733_),
    .B1(_13735_),
    .B2(_13626_),
    .ZN(_13736_));
 NOR4_X1 _23120_ (.A1(_13681_),
    .A2(_13729_),
    .A3(_13732_),
    .A4(_13736_),
    .ZN(_13737_));
 OR4_X1 _23121_ (.A1(_13714_),
    .A2(_13705_),
    .A3(_13727_),
    .A4(_13737_),
    .ZN(_00085_));
 NAND2_X1 _23122_ (.A1(_13353_),
    .A2(_13275_),
    .ZN(_13738_));
 AOI221_X2 _23123_ (.A(_13238_),
    .B1(_13275_),
    .B2(_13530_),
    .C1(_13738_),
    .C2(_13347_),
    .ZN(_13739_));
 AOI22_X1 _23124_ (.A1(_14987_),
    .A2(_13363_),
    .B1(_13720_),
    .B2(_14986_),
    .ZN(_13740_));
 OAI221_X1 _23125_ (.A(_13422_),
    .B1(_13723_),
    .B2(_14986_),
    .C1(_13740_),
    .C2(_15004_),
    .ZN(_13741_));
 OAI21_X1 _23126_ (.A(_13337_),
    .B1(_13275_),
    .B2(_13444_),
    .ZN(_13742_));
 AOI21_X1 _23127_ (.A(net141),
    .B1(_13585_),
    .B2(_13742_),
    .ZN(_13743_));
 AOI21_X1 _23128_ (.A(_13339_),
    .B1(_13667_),
    .B2(net141),
    .ZN(_13744_));
 OAI221_X2 _23129_ (.A(_13449_),
    .B1(_13744_),
    .B2(net175),
    .C1(net177),
    .C2(_13264_),
    .ZN(_13745_));
 AOI221_X2 _23130_ (.A(_13743_),
    .B1(_13720_),
    .B2(_13587_),
    .C1(_13363_),
    .C2(_13745_),
    .ZN(_13746_));
 OAI221_X1 _23131_ (.A(_13680_),
    .B1(_13739_),
    .B2(_13741_),
    .C1(_13746_),
    .C2(_13422_),
    .ZN(_13747_));
 NOR2_X1 _23132_ (.A1(_13228_),
    .A2(_13345_),
    .ZN(_13748_));
 NAND3_X1 _23133_ (.A1(_15011_),
    .A2(_13333_),
    .A3(_13604_),
    .ZN(_13749_));
 NAND3_X1 _23134_ (.A1(_13338_),
    .A2(_13283_),
    .A3(_13651_),
    .ZN(_13750_));
 AOI21_X1 _23135_ (.A(_13379_),
    .B1(_13749_),
    .B2(_13750_),
    .ZN(_13751_));
 OAI21_X1 _23136_ (.A(_13651_),
    .B1(_13257_),
    .B2(_14988_),
    .ZN(_13752_));
 AOI221_X1 _23137_ (.A(_13297_),
    .B1(_13752_),
    .B2(_13337_),
    .C1(_13278_),
    .C2(_13240_),
    .ZN(_13753_));
 NOR3_X1 _23138_ (.A1(_13371_),
    .A2(_13751_),
    .A3(_13753_),
    .ZN(_13754_));
 NOR2_X1 _23139_ (.A1(_15007_),
    .A2(_13495_),
    .ZN(_13755_));
 MUX2_X1 _23140_ (.A(_13353_),
    .B(_13350_),
    .S(_13217_),
    .Z(_13756_));
 AOI211_X2 _23141_ (.A(_13298_),
    .B(_13755_),
    .C1(_13756_),
    .C2(_13346_),
    .ZN(_13757_));
 AOI21_X1 _23142_ (.A(_13346_),
    .B1(_13512_),
    .B2(net178),
    .ZN(_13758_));
 NOR3_X1 _23143_ (.A1(_13380_),
    .A2(_13378_),
    .A3(_13758_),
    .ZN(_13759_));
 NOR3_X1 _23144_ (.A1(_13364_),
    .A2(_13757_),
    .A3(_13759_),
    .ZN(_13760_));
 OAI21_X1 _23145_ (.A(_13748_),
    .B1(_13754_),
    .B2(_13760_),
    .ZN(_13761_));
 AOI221_X2 _23146_ (.A(_13415_),
    .B1(_13287_),
    .B2(_13286_),
    .C1(net133),
    .C2(_13221_),
    .ZN(_13762_));
 NOR3_X1 _23147_ (.A1(_15005_),
    .A2(_15014_),
    .A3(_13334_),
    .ZN(_13763_));
 OAI21_X1 _23148_ (.A(_13379_),
    .B1(_13762_),
    .B2(_13763_),
    .ZN(_13764_));
 OR2_X1 _23149_ (.A1(_13337_),
    .A2(_13406_),
    .ZN(_13765_));
 OR2_X1 _23150_ (.A1(_13537_),
    .A2(_13444_),
    .ZN(_13766_));
 OAI221_X1 _23151_ (.A(_13298_),
    .B1(_13441_),
    .B2(_13765_),
    .C1(_13766_),
    .C2(_15011_),
    .ZN(_13767_));
 NAND3_X1 _23152_ (.A1(_13303_),
    .A2(_13764_),
    .A3(_13767_),
    .ZN(_13768_));
 NAND3_X1 _23153_ (.A1(_13238_),
    .A2(_13399_),
    .A3(_13372_),
    .ZN(_13769_));
 OAI221_X1 _23154_ (.A(_13223_),
    .B1(_13334_),
    .B2(_13603_),
    .C1(_13264_),
    .C2(net141),
    .ZN(_13770_));
 NAND3_X1 _23155_ (.A1(_13422_),
    .A2(_13769_),
    .A3(_13770_),
    .ZN(_13771_));
 OAI21_X1 _23156_ (.A(_13372_),
    .B1(_13346_),
    .B2(net177),
    .ZN(_13772_));
 OAI221_X1 _23157_ (.A(_13378_),
    .B1(_13442_),
    .B2(_13265_),
    .C1(_13772_),
    .C2(_15011_),
    .ZN(_13773_));
 NAND4_X1 _23158_ (.A1(_13236_),
    .A2(_13345_),
    .A3(_13771_),
    .A4(_13773_),
    .ZN(_13774_));
 AOI21_X1 _23159_ (.A(_13393_),
    .B1(_13238_),
    .B2(_13277_),
    .ZN(_13775_));
 AOI21_X1 _23160_ (.A(_13237_),
    .B1(_13411_),
    .B2(_13414_),
    .ZN(_13776_));
 NOR3_X1 _23161_ (.A1(_13463_),
    .A2(_13298_),
    .A3(_13776_),
    .ZN(_13777_));
 AOI21_X1 _23162_ (.A(_13638_),
    .B1(_13775_),
    .B2(_13777_),
    .ZN(_13778_));
 OAI221_X2 _23163_ (.A(_13614_),
    .B1(_13606_),
    .B2(_13338_),
    .C1(_13353_),
    .C2(_13328_),
    .ZN(_13779_));
 OAI221_X1 _23164_ (.A(_13493_),
    .B1(_13622_),
    .B2(_13530_),
    .C1(_13325_),
    .C2(_15011_),
    .ZN(_13780_));
 OR2_X1 _23165_ (.A1(_15006_),
    .A2(_13297_),
    .ZN(_13781_));
 OAI211_X2 _23166_ (.A(_13720_),
    .B(_13781_),
    .C1(_13378_),
    .C2(_13397_),
    .ZN(_13782_));
 NAND4_X1 _23167_ (.A1(_13778_),
    .A2(_13779_),
    .A3(_13780_),
    .A4(_13782_),
    .ZN(_13783_));
 AND3_X1 _23168_ (.A1(_13768_),
    .A2(_13774_),
    .A3(_13783_),
    .ZN(_13784_));
 NAND3_X1 _23169_ (.A1(_13747_),
    .A2(_13761_),
    .A3(_13784_),
    .ZN(_00086_));
 MUX2_X1 _23170_ (.A(net540),
    .B(_14992_),
    .S(_13218_),
    .Z(_13785_));
 OAI221_X1 _23171_ (.A(_13371_),
    .B1(_13734_),
    .B2(_13587_),
    .C1(_13785_),
    .C2(_13347_),
    .ZN(_13786_));
 AOI21_X1 _23172_ (.A(_13338_),
    .B1(_13283_),
    .B2(_13651_),
    .ZN(_13787_));
 OAI22_X1 _23173_ (.A1(net178),
    .A2(_13393_),
    .B1(_13604_),
    .B2(_13238_),
    .ZN(_13788_));
 OAI21_X1 _23174_ (.A(_13364_),
    .B1(_13787_),
    .B2(_13788_),
    .ZN(_13789_));
 NAND3_X1 _23175_ (.A1(_13363_),
    .A2(_13786_),
    .A3(_13789_),
    .ZN(_13790_));
 AOI21_X1 _23176_ (.A(_15004_),
    .B1(_13335_),
    .B2(_13340_),
    .ZN(_13791_));
 OR2_X1 _23177_ (.A1(_13371_),
    .A2(_13466_),
    .ZN(_13792_));
 NAND2_X1 _23178_ (.A1(_13240_),
    .A2(_13218_),
    .ZN(_13793_));
 MUX2_X1 _23179_ (.A(_15000_),
    .B(_13793_),
    .S(_13347_),
    .Z(_13794_));
 OAI221_X2 _23180_ (.A(_13345_),
    .B1(_13791_),
    .B2(_13792_),
    .C1(_13794_),
    .C2(_13364_),
    .ZN(_13795_));
 NAND3_X1 _23181_ (.A1(_13650_),
    .A2(_13790_),
    .A3(_13795_),
    .ZN(_13796_));
 AOI211_X2 _23182_ (.A(_13323_),
    .B(_13274_),
    .C1(_13481_),
    .C2(_13237_),
    .ZN(_13797_));
 OAI221_X2 _23183_ (.A(_13797_),
    .B1(_13328_),
    .B2(_13355_),
    .C1(_13353_),
    .C2(_13601_),
    .ZN(_13798_));
 NAND4_X1 _23184_ (.A1(net177),
    .A2(_14986_),
    .A3(_13362_),
    .A4(_13381_),
    .ZN(_13799_));
 AOI21_X1 _23185_ (.A(_13317_),
    .B1(_13334_),
    .B2(_13275_),
    .ZN(_13800_));
 OAI21_X1 _23186_ (.A(_13799_),
    .B1(_13800_),
    .B2(_13489_),
    .ZN(_13801_));
 OAI221_X2 _23187_ (.A(_13371_),
    .B1(_13463_),
    .B2(_13348_),
    .C1(_13383_),
    .C2(net611),
    .ZN(_13802_));
 OAI22_X1 _23188_ (.A1(_15011_),
    .A2(_13558_),
    .B1(_13654_),
    .B2(_13547_),
    .ZN(_13803_));
 OAI221_X2 _23189_ (.A(_13798_),
    .B1(_13801_),
    .B2(_13802_),
    .C1(_13803_),
    .C2(_13421_),
    .ZN(_13804_));
 MUX2_X1 _23190_ (.A(_13332_),
    .B(_13277_),
    .S(_13221_),
    .Z(_13805_));
 MUX2_X1 _23191_ (.A(_15014_),
    .B(_13805_),
    .S(_13495_),
    .Z(_13806_));
 OAI21_X1 _23192_ (.A(_13670_),
    .B1(_13654_),
    .B2(_13258_),
    .ZN(_13807_));
 MUX2_X1 _23193_ (.A(_13806_),
    .B(_13807_),
    .S(_13364_),
    .Z(_13808_));
 NOR2_X1 _23194_ (.A1(_13363_),
    .A2(_13404_),
    .ZN(_13809_));
 NOR2_X1 _23195_ (.A1(_13345_),
    .A2(_13404_),
    .ZN(_13810_));
 OAI21_X1 _23196_ (.A(_13464_),
    .B1(_13257_),
    .B2(_13177_),
    .ZN(_13811_));
 AOI21_X1 _23197_ (.A(_13435_),
    .B1(_13811_),
    .B2(_13348_),
    .ZN(_13812_));
 NOR2_X1 _23198_ (.A1(_13675_),
    .A2(_13762_),
    .ZN(_13813_));
 MUX2_X1 _23199_ (.A(_13812_),
    .B(_13813_),
    .S(_13235_),
    .Z(_13814_));
 AOI222_X2 _23200_ (.A1(_13562_),
    .A2(_13804_),
    .B1(_13809_),
    .B2(_13808_),
    .C1(_13810_),
    .C2(_13814_),
    .ZN(_13815_));
 AOI21_X1 _23201_ (.A(_13481_),
    .B1(_13278_),
    .B2(_14995_),
    .ZN(_13816_));
 OAI221_X1 _23202_ (.A(_13797_),
    .B1(_13816_),
    .B2(_14987_),
    .C1(_13328_),
    .C2(_13385_),
    .ZN(_13817_));
 OAI221_X1 _23203_ (.A(_13324_),
    .B1(_13674_),
    .B2(_15011_),
    .C1(_13382_),
    .C2(_13277_),
    .ZN(_13818_));
 AOI21_X1 _23204_ (.A(_13541_),
    .B1(_13817_),
    .B2(_13818_),
    .ZN(_13819_));
 NOR2_X1 _23205_ (.A1(_14987_),
    .A2(_13283_),
    .ZN(_13820_));
 AOI21_X1 _23206_ (.A(net178),
    .B1(_13288_),
    .B2(_13399_),
    .ZN(_13821_));
 OAI21_X1 _23207_ (.A(_13345_),
    .B1(_13820_),
    .B2(_13821_),
    .ZN(_13822_));
 AOI21_X1 _23208_ (.A(_13339_),
    .B1(_13381_),
    .B2(_14986_),
    .ZN(_13823_));
 NOR2_X1 _23209_ (.A1(_13278_),
    .A2(_13599_),
    .ZN(_13824_));
 OAI221_X1 _23210_ (.A(_13822_),
    .B1(_13823_),
    .B2(_13345_),
    .C1(_14987_),
    .C2(_13824_),
    .ZN(_13825_));
 NOR2_X1 _23211_ (.A1(_13364_),
    .A2(_13541_),
    .ZN(_13826_));
 AOI21_X1 _23212_ (.A(_13819_),
    .B1(_13825_),
    .B2(_13826_),
    .ZN(_13827_));
 NAND3_X1 _23213_ (.A1(_13815_),
    .A2(_13796_),
    .A3(_13827_),
    .ZN(_00087_));
 INV_X1 _23214_ (.A(net559),
    .ZN(_13828_));
 NOR2_X1 _23215_ (.A1(_13828_),
    .A2(_08994_),
    .ZN(_13829_));
 NOR2_X1 _23216_ (.A1(net559),
    .A2(_08994_),
    .ZN(_13830_));
 XNOR2_X2 _23217_ (.A(net657),
    .B(_11137_),
    .ZN(_13831_));
 XNOR2_X2 _23218_ (.A(_11183_),
    .B(_11120_),
    .ZN(_13832_));
 XNOR2_X2 _23219_ (.A(_13832_),
    .B(_11123_),
    .ZN(_13833_));
 XNOR2_X2 _23220_ (.A(_13833_),
    .B(_13831_),
    .ZN(_13834_));
 MUX2_X2 _23221_ (.A(_13829_),
    .B(_13830_),
    .S(_13834_),
    .Z(_13835_));
 NAND3_X1 _23222_ (.A1(net559),
    .A2(_09179_),
    .A3(_00461_),
    .ZN(_13836_));
 NAND2_X1 _23223_ (.A1(_13828_),
    .A2(_09728_),
    .ZN(_13837_));
 OAI21_X4 _23224_ (.A(_13836_),
    .B1(_13837_),
    .B2(_00461_),
    .ZN(_13838_));
 NOR2_X4 _23225_ (.A1(_13835_),
    .A2(_13838_),
    .ZN(_13839_));
 INV_X8 _23226_ (.A(net1186),
    .ZN(_13840_));
 BUF_X8 clone531 (.A(_14152_),
    .Z(net1115));
 BUF_X16 _23228_ (.A(_13840_),
    .Z(_15024_));
 XNOR2_X2 _23229_ (.A(_11135_),
    .B(\sa03_sr[0] ),
    .ZN(_13842_));
 XNOR2_X1 _23230_ (.A(_11136_),
    .B(net656),
    .ZN(_13843_));
 XOR2_X2 _23231_ (.A(_11120_),
    .B(_11183_),
    .Z(_13844_));
 NAND3_X1 _23232_ (.A1(net568),
    .A2(_09100_),
    .A3(_13844_),
    .ZN(_13845_));
 NOR2_X1 _23233_ (.A1(net568),
    .A2(_08993_),
    .ZN(_13846_));
 NAND2_X1 _23234_ (.A1(net970),
    .A2(_13846_),
    .ZN(_13847_));
 AOI21_X1 _23235_ (.A(_13843_),
    .B1(_13845_),
    .B2(_13847_),
    .ZN(_13848_));
 XOR2_X1 _23236_ (.A(_11136_),
    .B(net656),
    .Z(_13849_));
 NAND2_X1 _23237_ (.A1(_13844_),
    .A2(_13846_),
    .ZN(_13850_));
 NAND3_X1 _23238_ (.A1(net568),
    .A2(_09023_),
    .A3(net970),
    .ZN(_13851_));
 AOI21_X1 _23239_ (.A(_13849_),
    .B1(_13850_),
    .B2(_13851_),
    .ZN(_13852_));
 INV_X1 _23240_ (.A(net568),
    .ZN(_13853_));
 NAND3_X1 _23241_ (.A1(_13853_),
    .A2(_09030_),
    .A3(_00462_),
    .ZN(_13854_));
 NAND2_X1 _23242_ (.A1(net568),
    .A2(_09102_),
    .ZN(_13855_));
 OAI21_X1 _23243_ (.A(_13854_),
    .B1(_13855_),
    .B2(_00462_),
    .ZN(_13856_));
 OR3_X4 _23244_ (.A1(_13848_),
    .A2(_13852_),
    .A3(_13856_),
    .ZN(_13857_));
 INV_X8 _23245_ (.A(_13857_),
    .ZN(_13858_));
 BUF_X8 _23246_ (.A(_13858_),
    .Z(_13859_));
 BUF_X8 _23247_ (.A(_13859_),
    .Z(_15027_));
 XOR2_X2 _23248_ (.A(_11114_),
    .B(_11159_),
    .Z(_13860_));
 XOR2_X2 _23249_ (.A(net972),
    .B(_13860_),
    .Z(_13861_));
 XOR2_X2 _23250_ (.A(_11164_),
    .B(_11219_),
    .Z(_13862_));
 NAND3_X1 _23251_ (.A1(_06295_),
    .A2(net949),
    .A3(_13862_),
    .ZN(_13863_));
 XNOR2_X2 _23252_ (.A(_11164_),
    .B(_11219_),
    .ZN(_13864_));
 NOR2_X1 _23253_ (.A1(_06295_),
    .A2(_09015_),
    .ZN(_13865_));
 NAND2_X1 _23254_ (.A1(_13864_),
    .A2(_13865_),
    .ZN(_13866_));
 AOI21_X2 _23255_ (.A(_13861_),
    .B1(_13863_),
    .B2(_13866_),
    .ZN(_13867_));
 XNOR2_X1 _23256_ (.A(net972),
    .B(_13860_),
    .ZN(_13868_));
 NAND2_X1 _23257_ (.A1(_13862_),
    .A2(_13865_),
    .ZN(_13869_));
 NAND3_X1 _23258_ (.A1(_06295_),
    .A2(_09194_),
    .A3(_13864_),
    .ZN(_13870_));
 AOI21_X2 _23259_ (.A(_13868_),
    .B1(_13869_),
    .B2(_13870_),
    .ZN(_13871_));
 NAND3_X1 _23260_ (.A1(_06308_),
    .A2(_09727_),
    .A3(_00463_),
    .ZN(_13872_));
 NAND2_X1 _23261_ (.A1(_06295_),
    .A2(_09028_),
    .ZN(_13873_));
 OAI21_X2 _23262_ (.A(_13872_),
    .B1(_13873_),
    .B2(_00463_),
    .ZN(_13874_));
 NOR3_X4 _23263_ (.A1(_13867_),
    .A2(_13871_),
    .A3(_13874_),
    .ZN(_13875_));
 INV_X4 _23264_ (.A(_13875_),
    .ZN(_13876_));
 BUF_X4 _23265_ (.A(_13876_),
    .Z(_13877_));
 BUF_X4 _23266_ (.A(_13877_),
    .Z(_13878_));
 BUF_X4 _23267_ (.A(_13878_),
    .Z(_13879_));
 BUF_X4 _23268_ (.A(_13879_),
    .Z(_15043_));
 BUF_X8 _23269_ (.A(_13857_),
    .Z(_13880_));
 BUF_X8 _23270_ (.A(_13880_),
    .Z(_15018_));
 BUF_X4 _23271_ (.A(net962),
    .Z(_13881_));
 BUF_X4 _23272_ (.A(_13881_),
    .Z(_13882_));
 BUF_X4 _23273_ (.A(_13882_),
    .Z(_13883_));
 BUF_X4 _23274_ (.A(_13883_),
    .Z(_15036_));
 INV_X1 _23275_ (.A(_06268_),
    .ZN(_13884_));
 XNOR2_X1 _23276_ (.A(_11246_),
    .B(_11202_),
    .ZN(_13885_));
 NOR3_X1 _23277_ (.A1(_13884_),
    .A2(_09823_),
    .A3(_13885_),
    .ZN(_13886_));
 NOR3_X1 _23278_ (.A1(_06268_),
    .A2(_09823_),
    .A3(_13885_),
    .ZN(_13887_));
 MUX2_X2 _23279_ (.A(_13886_),
    .B(_13887_),
    .S(_11264_),
    .Z(_13888_));
 XOR2_X2 _23280_ (.A(_11246_),
    .B(_11202_),
    .Z(_13889_));
 NOR3_X1 _23281_ (.A1(_06268_),
    .A2(_08975_),
    .A3(_13889_),
    .ZN(_13890_));
 NOR3_X1 _23282_ (.A1(_13884_),
    .A2(_08975_),
    .A3(_13889_),
    .ZN(_13891_));
 MUX2_X1 _23283_ (.A(_13890_),
    .B(_13891_),
    .S(_11264_),
    .Z(_13892_));
 NAND3_X1 _23284_ (.A1(_06268_),
    .A2(_08996_),
    .A3(\text_in_r[21] ),
    .ZN(_13893_));
 NAND2_X1 _23285_ (.A1(_13884_),
    .A2(_08996_),
    .ZN(_13894_));
 OAI21_X2 _23286_ (.A(_13893_),
    .B1(_13894_),
    .B2(\text_in_r[21] ),
    .ZN(_13895_));
 OR3_X2 _23287_ (.A1(_13888_),
    .A2(_13892_),
    .A3(_13895_),
    .ZN(_13896_));
 BUF_X4 _23288_ (.A(_13896_),
    .Z(_13897_));
 CLKBUF_X3 _23289_ (.A(_13897_),
    .Z(_13898_));
 XNOR2_X1 _23290_ (.A(_11185_),
    .B(_11200_),
    .ZN(_13899_));
 XNOR2_X1 _23291_ (.A(_11119_),
    .B(_13899_),
    .ZN(_13900_));
 MUX2_X2 _23292_ (.A(\text_in_r[23] ),
    .B(_13900_),
    .S(_09803_),
    .Z(_13901_));
 XOR2_X2 _23293_ (.A(_06586_),
    .B(_13901_),
    .Z(_13902_));
 XNOR2_X1 _23294_ (.A(_11201_),
    .B(_11199_),
    .ZN(_13903_));
 XNOR2_X2 _23295_ (.A(_11198_),
    .B(_11187_),
    .ZN(_13904_));
 XNOR2_X1 _23296_ (.A(_11261_),
    .B(_13904_),
    .ZN(_13905_));
 XNOR2_X1 _23297_ (.A(_13903_),
    .B(_13905_),
    .ZN(_13906_));
 MUX2_X2 _23298_ (.A(\text_in_r[22] ),
    .B(_13906_),
    .S(_11207_),
    .Z(_13907_));
 XNOR2_X2 _23299_ (.A(_06574_),
    .B(_13907_),
    .ZN(_13908_));
 BUF_X4 _23300_ (.A(_13908_),
    .Z(_13909_));
 INV_X1 _23301_ (.A(_06285_),
    .ZN(_13910_));
 NOR2_X1 _23302_ (.A1(_13910_),
    .A2(_09823_),
    .ZN(_13911_));
 NOR2_X1 _23303_ (.A1(_06285_),
    .A2(_09823_),
    .ZN(_13912_));
 XNOR2_X1 _23304_ (.A(_11250_),
    .B(_11183_),
    .ZN(_13913_));
 XNOR2_X1 _23305_ (.A(_11220_),
    .B(_13913_),
    .ZN(_13914_));
 XOR2_X1 _23306_ (.A(_11246_),
    .B(_11265_),
    .Z(_13915_));
 XNOR2_X1 _23307_ (.A(_11224_),
    .B(_13915_),
    .ZN(_13916_));
 XNOR2_X1 _23308_ (.A(_13914_),
    .B(_13916_),
    .ZN(_13917_));
 MUX2_X2 _23309_ (.A(_13911_),
    .B(_13912_),
    .S(_13917_),
    .Z(_13918_));
 NAND3_X2 _23310_ (.A1(_13910_),
    .A2(_09135_),
    .A3(\text_in_r[20] ),
    .ZN(_13919_));
 NAND2_X1 _23311_ (.A1(_06285_),
    .A2(_09180_),
    .ZN(_13920_));
 OAI21_X4 _23312_ (.A(_13919_),
    .B1(_13920_),
    .B2(\text_in_r[20] ),
    .ZN(_13921_));
 NOR2_X4 _23313_ (.A1(_13918_),
    .A2(_13921_),
    .ZN(_13922_));
 BUF_X4 _23314_ (.A(_13922_),
    .Z(_13923_));
 BUF_X4 _23315_ (.A(_13923_),
    .Z(_13924_));
 NOR2_X1 _23316_ (.A1(_13909_),
    .A2(_13924_),
    .ZN(_13925_));
 BUF_X4 _23317_ (.A(_15021_),
    .Z(_13926_));
 NAND2_X1 _23318_ (.A1(_06229_),
    .A2(_11191_),
    .ZN(_13927_));
 INV_X1 _23319_ (.A(_06229_),
    .ZN(_13928_));
 NAND2_X1 _23320_ (.A1(_13928_),
    .A2(_09076_),
    .ZN(_13929_));
 XNOR2_X2 _23321_ (.A(_11159_),
    .B(_11225_),
    .ZN(_13930_));
 XNOR2_X1 _23322_ (.A(_13844_),
    .B(_13930_),
    .ZN(_13931_));
 XOR2_X1 _23323_ (.A(_11220_),
    .B(_11245_),
    .Z(_13932_));
 XNOR2_X1 _23324_ (.A(_11158_),
    .B(_13932_),
    .ZN(_13933_));
 XNOR2_X2 _23325_ (.A(_13931_),
    .B(_13933_),
    .ZN(_13934_));
 MUX2_X2 _23326_ (.A(_13927_),
    .B(_13929_),
    .S(_13934_),
    .Z(_13935_));
 CLKBUF_X3 _23327_ (.A(\text_in_r[19] ),
    .Z(_13936_));
 NAND2_X2 _23328_ (.A1(_06229_),
    .A2(net610),
    .ZN(_13937_));
 NOR2_X1 _23329_ (.A1(_13936_),
    .A2(_13937_),
    .ZN(_13938_));
 NOR2_X2 _23330_ (.A1(_06229_),
    .A2(net594),
    .ZN(_13939_));
 AOI21_X4 _23331_ (.A(_13938_),
    .B1(_13939_),
    .B2(_13936_),
    .ZN(_13940_));
 AOI21_X4 _23332_ (.A(_13926_),
    .B1(_13935_),
    .B2(_13940_),
    .ZN(_13941_));
 NOR2_X1 _23333_ (.A1(_13928_),
    .A2(_08974_),
    .ZN(_13942_));
 NOR2_X1 _23334_ (.A1(_06229_),
    .A2(_08974_),
    .ZN(_13943_));
 MUX2_X2 _23335_ (.A(_13942_),
    .B(_13943_),
    .S(_13934_),
    .Z(_13944_));
 BUF_X8 _23336_ (.A(_13944_),
    .Z(_13945_));
 NAND2_X1 _23337_ (.A1(_13936_),
    .A2(_13939_),
    .ZN(_13946_));
 OAI21_X4 _23338_ (.A(_13946_),
    .B1(_13937_),
    .B2(_13936_),
    .ZN(_13947_));
 BUF_X8 _23339_ (.A(_13947_),
    .Z(_13948_));
 NOR2_X4 _23340_ (.A1(_13945_),
    .A2(_13948_),
    .ZN(_13949_));
 BUF_X4 _23341_ (.A(_13949_),
    .Z(_13950_));
 BUF_X4 _23342_ (.A(_13950_),
    .Z(_13951_));
 BUF_X4 _23343_ (.A(_15030_),
    .Z(_13952_));
 INV_X2 _23344_ (.A(_13952_),
    .ZN(_13953_));
 AOI21_X1 _23345_ (.A(_13941_),
    .B1(_13951_),
    .B2(_13953_),
    .ZN(_13954_));
 BUF_X2 clone187 (.A(_15204_),
    .Z(net187));
 BUF_X4 _23347_ (.A(net967),
    .Z(_13956_));
 BUF_X8 _23348_ (.A(_13935_),
    .Z(_13957_));
 BUF_X8 _23349_ (.A(_13940_),
    .Z(_13958_));
 NAND3_X1 _23350_ (.A1(_13876_),
    .A2(_13957_),
    .A3(_13958_),
    .ZN(_13959_));
 BUF_X4 _23351_ (.A(_13959_),
    .Z(_13960_));
 OAI221_X1 _23352_ (.A(_13925_),
    .B1(_13954_),
    .B2(_13879_),
    .C1(_13956_),
    .C2(_13960_),
    .ZN(_13961_));
 OR2_X1 _23353_ (.A1(_13918_),
    .A2(_13921_),
    .ZN(_13962_));
 CLKBUF_X3 _23354_ (.A(_13962_),
    .Z(_13963_));
 BUF_X4 _23355_ (.A(_13963_),
    .Z(_13964_));
 BUF_X4 _23356_ (.A(_13877_),
    .Z(_13965_));
 NAND2_X4 _23357_ (.A1(_13935_),
    .A2(_13940_),
    .ZN(_13966_));
 BUF_X4 _23358_ (.A(_13966_),
    .Z(_13967_));
 OAI21_X4 _23359_ (.A(_13859_),
    .B1(_13838_),
    .B2(net958),
    .ZN(_13968_));
 AOI21_X1 _23360_ (.A(_13965_),
    .B1(_13967_),
    .B2(_13968_),
    .ZN(_13969_));
 BUF_X4 _23361_ (.A(_13945_),
    .Z(_13970_));
 BUF_X4 _23362_ (.A(_13948_),
    .Z(_13971_));
 OAI21_X4 _23363_ (.A(_13876_),
    .B1(_13970_),
    .B2(_13971_),
    .ZN(_13972_));
 OAI22_X2 _23364_ (.A1(_13956_),
    .A2(_13967_),
    .B1(_13972_),
    .B2(_13859_),
    .ZN(_13973_));
 NOR3_X1 _23365_ (.A1(_13964_),
    .A2(_13969_),
    .A3(_13973_),
    .ZN(_13974_));
 NAND3_X1 _23366_ (.A1(_15022_),
    .A2(_13935_),
    .A3(_13940_),
    .ZN(_13975_));
 OAI21_X4 _23367_ (.A(_13858_),
    .B1(_13945_),
    .B2(_13948_),
    .ZN(_13976_));
 AND2_X1 _23368_ (.A1(_13975_),
    .A2(_13976_),
    .ZN(_13977_));
 AOI21_X1 _23369_ (.A(net964),
    .B1(_13949_),
    .B2(net967),
    .ZN(_13978_));
 NOR2_X2 clone149 (.A1(_13838_),
    .A2(_13835_),
    .ZN(net149));
 INV_X2 _23371_ (.A(_15020_),
    .ZN(_13980_));
 NAND3_X4 _23372_ (.A1(_13857_),
    .A2(_13957_),
    .A3(_13958_),
    .ZN(_13981_));
 OAI22_X1 _23373_ (.A1(_13980_),
    .A2(_13949_),
    .B1(_13981_),
    .B2(net149),
    .ZN(_13982_));
 AOI221_X2 _23374_ (.A(_13963_),
    .B1(_13977_),
    .B2(_13978_),
    .C1(_13982_),
    .C2(_13882_),
    .ZN(_13983_));
 NOR3_X4 _23375_ (.A1(_13875_),
    .A2(_13945_),
    .A3(_13948_),
    .ZN(_13984_));
 BUF_X16 _23376_ (.A(net969),
    .Z(_13985_));
 AOI22_X1 _23377_ (.A1(_15041_),
    .A2(_13967_),
    .B1(_13984_),
    .B2(_13985_),
    .ZN(_13986_));
 OAI21_X1 _23378_ (.A(_13908_),
    .B1(_13924_),
    .B2(_13986_),
    .ZN(_13987_));
 OAI22_X1 _23379_ (.A1(_13909_),
    .A2(_13974_),
    .B1(_13983_),
    .B2(_13987_),
    .ZN(_13988_));
 AND4_X1 _23380_ (.A1(_13898_),
    .A2(_13902_),
    .A3(_13961_),
    .A4(_13988_),
    .ZN(_13989_));
 NOR3_X4 _23381_ (.A1(_13888_),
    .A2(_13892_),
    .A3(_13895_),
    .ZN(_13990_));
 BUF_X4 _23382_ (.A(_13990_),
    .Z(_13991_));
 BUF_X4 _23383_ (.A(_13991_),
    .Z(_13992_));
 CLKBUF_X3 _23384_ (.A(_13902_),
    .Z(_13993_));
 XOR2_X2 _23385_ (.A(_06574_),
    .B(_13907_),
    .Z(_13994_));
 INV_X8 _23386_ (.A(_13926_),
    .ZN(_13995_));
 NOR3_X4 _23387_ (.A1(_13995_),
    .A2(_13945_),
    .A3(_13948_),
    .ZN(_13996_));
 NAND2_X1 _23388_ (.A1(_13839_),
    .A2(_13876_),
    .ZN(_13997_));
 NOR2_X2 _23389_ (.A1(net969),
    .A2(net964),
    .ZN(_13998_));
 NAND2_X2 _23390_ (.A1(net149),
    .A2(_13949_),
    .ZN(_13999_));
 AOI221_X2 _23391_ (.A(_13922_),
    .B1(_13996_),
    .B2(_13997_),
    .C1(_13998_),
    .C2(_13999_),
    .ZN(_14000_));
 BUF_X4 _23392_ (.A(_15028_),
    .Z(_14001_));
 NAND2_X1 _23393_ (.A1(_14001_),
    .A2(_13984_),
    .ZN(_14002_));
 AOI21_X4 _23394_ (.A(net963),
    .B1(_13935_),
    .B2(_13940_),
    .ZN(_14003_));
 NOR3_X4 _23395_ (.A1(_13876_),
    .A2(_13945_),
    .A3(_13948_),
    .ZN(_14004_));
 NOR2_X4 _23396_ (.A1(_14003_),
    .A2(_14004_),
    .ZN(_14005_));
 OAI21_X4 _23397_ (.A(_13881_),
    .B1(_13970_),
    .B2(_13971_),
    .ZN(_14006_));
 OAI221_X2 _23398_ (.A(_14002_),
    .B1(_14005_),
    .B2(_13980_),
    .C1(_14006_),
    .C2(_13985_),
    .ZN(_14007_));
 AOI211_X2 _23399_ (.A(_13994_),
    .B(_14000_),
    .C1(_14007_),
    .C2(_13924_),
    .ZN(_14008_));
 NOR3_X1 _23400_ (.A1(_13992_),
    .A2(_13993_),
    .A3(_14008_),
    .ZN(_14009_));
 CLKBUF_X3 _23401_ (.A(_13994_),
    .Z(_14010_));
 BUF_X4 _23402_ (.A(_13963_),
    .Z(_14011_));
 BUF_X4 _23403_ (.A(_14011_),
    .Z(_14012_));
 NAND2_X1 _23404_ (.A1(_13880_),
    .A2(_13965_),
    .ZN(_14013_));
 BUF_X4 _23405_ (.A(_13840_),
    .Z(_14014_));
 CLKBUF_X3 _23406_ (.A(_13967_),
    .Z(_14015_));
 NOR2_X1 _23407_ (.A1(_14014_),
    .A2(_14015_),
    .ZN(_14016_));
 BUF_X8 _23408_ (.A(_15034_),
    .Z(_14017_));
 BUF_X4 _23409_ (.A(_13949_),
    .Z(_14018_));
 MUX2_X1 _23410_ (.A(_14017_),
    .B(_14014_),
    .S(_14018_),
    .Z(_14019_));
 BUF_X4 _23411_ (.A(_13876_),
    .Z(_14020_));
 BUF_X4 _23412_ (.A(_14020_),
    .Z(_14021_));
 BUF_X4 _23413_ (.A(_14021_),
    .Z(_14022_));
 OAI221_X2 _23414_ (.A(_14012_),
    .B1(_14013_),
    .B2(_14016_),
    .C1(_14019_),
    .C2(_14022_),
    .ZN(_14023_));
 BUF_X8 _23415_ (.A(_15022_),
    .Z(_14024_));
 NAND2_X1 _23416_ (.A1(_13883_),
    .A2(_13951_),
    .ZN(_14025_));
 NOR2_X4 _23417_ (.A1(_13857_),
    .A2(_13876_),
    .ZN(_14026_));
 AOI21_X1 _23418_ (.A(_13984_),
    .B1(_14026_),
    .B2(_14015_),
    .ZN(_14027_));
 BUF_X4 _23419_ (.A(_13839_),
    .Z(_14028_));
 BUF_X4 _23420_ (.A(_14028_),
    .Z(_14029_));
 OAI222_X2 _23421_ (.A1(_14024_),
    .A2(_14025_),
    .B1(_14027_),
    .B2(_14029_),
    .C1(_15027_),
    .C2(_13972_),
    .ZN(_14030_));
 BUF_X4 _23422_ (.A(_13964_),
    .Z(_14031_));
 OAI21_X1 _23423_ (.A(_14023_),
    .B1(_14030_),
    .B2(_14031_),
    .ZN(_14032_));
 NAND2_X1 _23424_ (.A1(_14010_),
    .A2(_14032_),
    .ZN(_14033_));
 BUF_X4 _23425_ (.A(_13897_),
    .Z(_14034_));
 NOR2_X1 _23426_ (.A1(_14034_),
    .A2(_13902_),
    .ZN(_14035_));
 BUF_X4 _23427_ (.A(_13966_),
    .Z(_14036_));
 OAI221_X1 _23428_ (.A(_14011_),
    .B1(_14006_),
    .B2(_13995_),
    .C1(_13880_),
    .C2(_14036_),
    .ZN(_14037_));
 AOI21_X4 _23429_ (.A(_14017_),
    .B1(_13957_),
    .B2(_13958_),
    .ZN(_14038_));
 CLKBUF_X3 _23430_ (.A(_14018_),
    .Z(_14039_));
 AOI21_X1 _23431_ (.A(_14038_),
    .B1(_14039_),
    .B2(_14014_),
    .ZN(_14040_));
 AOI21_X1 _23432_ (.A(_14037_),
    .B1(_14040_),
    .B2(_14022_),
    .ZN(_14041_));
 NOR2_X2 _23433_ (.A1(_14014_),
    .A2(_14018_),
    .ZN(_14042_));
 NOR3_X2 _23434_ (.A1(_13859_),
    .A2(_13918_),
    .A3(_13921_),
    .ZN(_14043_));
 NAND2_X1 _23435_ (.A1(_13878_),
    .A2(_14043_),
    .ZN(_14044_));
 NAND2_X2 _23436_ (.A1(_13967_),
    .A2(_13922_),
    .ZN(_14045_));
 INV_X4 _23437_ (.A(net968),
    .ZN(_14046_));
 BUF_X4 _23438_ (.A(_13881_),
    .Z(_14047_));
 NAND2_X1 _23439_ (.A1(_14046_),
    .A2(_14047_),
    .ZN(_14048_));
 OAI221_X2 _23440_ (.A(_13994_),
    .B1(_14042_),
    .B2(_14044_),
    .C1(_14045_),
    .C2(_14048_),
    .ZN(_14049_));
 OAI21_X1 _23441_ (.A(_14035_),
    .B1(_14041_),
    .B2(_14049_),
    .ZN(_14050_));
 BUF_X4 _23442_ (.A(_13923_),
    .Z(_14051_));
 NAND2_X1 _23443_ (.A1(net572),
    .A2(_13984_),
    .ZN(_14052_));
 NOR3_X4 _23444_ (.A1(net1207),
    .A2(_13945_),
    .A3(_13948_),
    .ZN(_14053_));
 AOI21_X4 _23445_ (.A(net968),
    .B1(_13957_),
    .B2(_13958_),
    .ZN(_14054_));
 OAI21_X1 _23446_ (.A(_15036_),
    .B1(_14053_),
    .B2(_14054_),
    .ZN(_14055_));
 AOI21_X1 _23447_ (.A(_14051_),
    .B1(_14052_),
    .B2(_14055_),
    .ZN(_14056_));
 OAI21_X2 _23448_ (.A(_13875_),
    .B1(_13838_),
    .B2(_13835_),
    .ZN(_14057_));
 AOI21_X4 _23449_ (.A(_13966_),
    .B1(_13877_),
    .B2(_13985_),
    .ZN(_14058_));
 NAND2_X4 _23450_ (.A1(_13859_),
    .A2(net965),
    .ZN(_14059_));
 OAI21_X1 _23451_ (.A(_14059_),
    .B1(_14047_),
    .B2(_14001_),
    .ZN(_14060_));
 BUF_X4 _23452_ (.A(_13967_),
    .Z(_14061_));
 AOI221_X2 _23453_ (.A(_14011_),
    .B1(_14057_),
    .B2(_14058_),
    .C1(_14060_),
    .C2(_14061_),
    .ZN(_14062_));
 NOR2_X1 _23454_ (.A1(_14056_),
    .A2(_14062_),
    .ZN(_14063_));
 NAND3_X1 _23455_ (.A1(_14010_),
    .A2(_14050_),
    .A3(_14063_),
    .ZN(_14064_));
 BUF_X4 _23456_ (.A(_13990_),
    .Z(_14065_));
 NAND2_X2 _23457_ (.A1(_14065_),
    .A2(_13902_),
    .ZN(_14066_));
 NOR3_X2 _23458_ (.A1(_13859_),
    .A2(_13945_),
    .A3(_13948_),
    .ZN(_14067_));
 NAND2_X2 _23459_ (.A1(_13840_),
    .A2(_14067_),
    .ZN(_14068_));
 INV_X2 _23460_ (.A(_14024_),
    .ZN(_14069_));
 AOI21_X4 _23461_ (.A(_13877_),
    .B1(_13966_),
    .B2(_14069_),
    .ZN(_14070_));
 INV_X1 _23462_ (.A(_14001_),
    .ZN(_14071_));
 AOI221_X1 _23463_ (.A(_13923_),
    .B1(_14068_),
    .B2(_14070_),
    .C1(_13984_),
    .C2(_14071_),
    .ZN(_14072_));
 AOI21_X4 _23464_ (.A(_13858_),
    .B1(_13935_),
    .B2(_13940_),
    .ZN(_14073_));
 NAND2_X4 _23465_ (.A1(net1185),
    .A2(_14073_),
    .ZN(_14074_));
 NOR2_X1 _23466_ (.A1(_14020_),
    .A2(_14053_),
    .ZN(_14075_));
 AOI221_X1 _23467_ (.A(_14011_),
    .B1(_14074_),
    .B2(_14075_),
    .C1(_14003_),
    .C2(_13952_),
    .ZN(_14076_));
 NOR3_X1 _23468_ (.A1(_13994_),
    .A2(_14072_),
    .A3(_14076_),
    .ZN(_14077_));
 NOR3_X4 _23469_ (.A1(_13857_),
    .A2(_13944_),
    .A3(_13947_),
    .ZN(_14078_));
 NAND2_X1 _23470_ (.A1(_13840_),
    .A2(_14078_),
    .ZN(_14079_));
 AOI21_X1 _23471_ (.A(net964),
    .B1(_13966_),
    .B2(_15020_),
    .ZN(_14080_));
 NOR3_X4 _23472_ (.A1(_13926_),
    .A2(_13945_),
    .A3(_13948_),
    .ZN(_14081_));
 AOI21_X1 _23473_ (.A(_14081_),
    .B1(_13966_),
    .B2(_15028_),
    .ZN(_14082_));
 AOI221_X2 _23474_ (.A(_13963_),
    .B1(_14079_),
    .B2(_14080_),
    .C1(_14082_),
    .C2(_13881_),
    .ZN(_14083_));
 AOI21_X1 _23475_ (.A(_14026_),
    .B1(_13880_),
    .B2(net149),
    .ZN(_14084_));
 XNOR2_X1 _23476_ (.A(_14036_),
    .B(_14084_),
    .ZN(_14085_));
 AOI211_X2 _23477_ (.A(_13994_),
    .B(_14083_),
    .C1(_14085_),
    .C2(_13964_),
    .ZN(_14086_));
 OAI22_X2 _23478_ (.A1(_14066_),
    .A2(_14077_),
    .B1(_14086_),
    .B2(_14050_),
    .ZN(_14087_));
 AOI221_X2 _23479_ (.A(_13989_),
    .B1(_14009_),
    .B2(_14033_),
    .C1(_14064_),
    .C2(_14087_),
    .ZN(_00088_));
 BUF_X4 _23480_ (.A(_14031_),
    .Z(_14088_));
 BUF_X4 _23481_ (.A(_14078_),
    .Z(_14089_));
 NOR3_X1 _23482_ (.A1(_13878_),
    .A2(_14089_),
    .A3(_14054_),
    .ZN(_14090_));
 XNOR2_X2 _23483_ (.A(net961),
    .B(_13950_),
    .ZN(_14091_));
 AOI21_X1 _23484_ (.A(_14090_),
    .B1(_14091_),
    .B2(_15043_),
    .ZN(_14092_));
 NOR2_X2 _23485_ (.A1(_14028_),
    .A2(_14018_),
    .ZN(_14093_));
 NOR2_X1 _23486_ (.A1(_13880_),
    .A2(_13882_),
    .ZN(_14094_));
 NOR2_X2 _23487_ (.A1(_13859_),
    .A2(_13876_),
    .ZN(_14095_));
 NOR2_X1 _23488_ (.A1(_14094_),
    .A2(_14095_),
    .ZN(_14096_));
 AND2_X1 _23489_ (.A1(_14093_),
    .A2(_14096_),
    .ZN(_14097_));
 CLKBUF_X3 _23490_ (.A(_14061_),
    .Z(_14098_));
 NAND2_X2 _23491_ (.A1(_13880_),
    .A2(_13881_),
    .ZN(_14099_));
 NAND2_X1 _23492_ (.A1(net571),
    .A2(_13877_),
    .ZN(_14100_));
 AOI21_X1 _23493_ (.A(_14098_),
    .B1(_14099_),
    .B2(_14100_),
    .ZN(_14101_));
 OR2_X1 _23494_ (.A1(_13898_),
    .A2(_14101_),
    .ZN(_14102_));
 OAI221_X1 _23495_ (.A(_14088_),
    .B1(_13992_),
    .B2(_14092_),
    .C1(_14097_),
    .C2(_14102_),
    .ZN(_14103_));
 XNOR2_X2 _23496_ (.A(_06586_),
    .B(_13901_),
    .ZN(_14104_));
 NAND2_X2 _23497_ (.A1(_13909_),
    .A2(_14104_),
    .ZN(_14105_));
 MUX2_X1 _23498_ (.A(_14071_),
    .B(_13968_),
    .S(_13881_),
    .Z(_14106_));
 AOI21_X1 _23499_ (.A(_13964_),
    .B1(_14106_),
    .B2(_14039_),
    .ZN(_14107_));
 CLKBUF_X3 _23500_ (.A(_13951_),
    .Z(_14108_));
 OR3_X1 _23501_ (.A1(_15044_),
    .A2(_14108_),
    .A3(_13991_),
    .ZN(_14109_));
 AOI21_X1 _23502_ (.A(_14105_),
    .B1(_14107_),
    .B2(_14109_),
    .ZN(_14110_));
 AOI21_X4 _23503_ (.A(_13995_),
    .B1(_13957_),
    .B2(_13958_),
    .ZN(_14111_));
 OAI21_X2 _23504_ (.A(_13878_),
    .B1(_14089_),
    .B2(_14111_),
    .ZN(_14112_));
 AOI21_X4 _23505_ (.A(_13876_),
    .B1(_13957_),
    .B2(_13958_),
    .ZN(_14113_));
 NAND2_X1 _23506_ (.A1(_13980_),
    .A2(_14113_),
    .ZN(_14114_));
 AND3_X1 _23507_ (.A1(_13991_),
    .A2(_14112_),
    .A3(_14114_),
    .ZN(_14115_));
 AND2_X1 _23508_ (.A1(_14003_),
    .A2(_13968_),
    .ZN(_14116_));
 INV_X2 _23509_ (.A(_15034_),
    .ZN(_14117_));
 AOI21_X1 _23510_ (.A(_13975_),
    .B1(_13883_),
    .B2(_14117_),
    .ZN(_14118_));
 BUF_X4 _23511_ (.A(_13965_),
    .Z(_14119_));
 OAI21_X4 _23512_ (.A(_13995_),
    .B1(_13970_),
    .B2(_13971_),
    .ZN(_14120_));
 NAND3_X2 _23513_ (.A1(_14017_),
    .A2(_13957_),
    .A3(_13958_),
    .ZN(_14121_));
 AOI21_X2 _23514_ (.A(_14119_),
    .B1(_14120_),
    .B2(_14121_),
    .ZN(_14122_));
 NOR4_X4 _23515_ (.A1(_14116_),
    .A2(_14122_),
    .A3(_14118_),
    .A4(_13992_),
    .ZN(_14123_));
 OAI21_X1 _23516_ (.A(_14004_),
    .B1(_13992_),
    .B2(net1183),
    .ZN(_14124_));
 OAI221_X2 _23517_ (.A(_14088_),
    .B1(_14123_),
    .B2(_14115_),
    .C1(_14124_),
    .C2(_14069_),
    .ZN(_14125_));
 NAND2_X2 _23518_ (.A1(_13994_),
    .A2(_14104_),
    .ZN(_14126_));
 NOR3_X2 _23519_ (.A1(net570),
    .A2(_13970_),
    .A3(_13971_),
    .ZN(_14127_));
 OAI21_X1 _23520_ (.A(_13879_),
    .B1(_14093_),
    .B2(_14127_),
    .ZN(_14128_));
 OR3_X4 _23521_ (.A1(_13918_),
    .A2(_13921_),
    .A3(_13896_),
    .ZN(_14129_));
 NOR2_X1 _23522_ (.A1(_14090_),
    .A2(_14129_),
    .ZN(_14130_));
 AOI21_X1 _23523_ (.A(_13941_),
    .B1(_14089_),
    .B2(_14014_),
    .ZN(_14131_));
 OAI22_X1 _23524_ (.A1(_15027_),
    .A2(_13960_),
    .B1(_14131_),
    .B2(_14022_),
    .ZN(_14132_));
 NOR2_X2 _23525_ (.A1(_14011_),
    .A2(_13990_),
    .ZN(_14133_));
 AOI221_X1 _23526_ (.A(_14126_),
    .B1(_14128_),
    .B2(_14130_),
    .C1(_14132_),
    .C2(_14133_),
    .ZN(_14134_));
 AOI22_X2 _23527_ (.A1(_14103_),
    .A2(_14110_),
    .B1(_14125_),
    .B2(_14134_),
    .ZN(_14135_));
 NAND2_X1 _23528_ (.A1(_14031_),
    .A2(_14034_),
    .ZN(_14136_));
 AOI21_X4 _23529_ (.A(_14046_),
    .B1(_13957_),
    .B2(_13958_),
    .ZN(_14137_));
 NOR3_X1 _23530_ (.A1(_15036_),
    .A2(_14089_),
    .A3(_14137_),
    .ZN(_14138_));
 NOR3_X1 _23531_ (.A1(_14022_),
    .A2(_13941_),
    .A3(_14127_),
    .ZN(_14139_));
 NOR3_X1 _23532_ (.A1(_14136_),
    .A2(_14138_),
    .A3(_14139_),
    .ZN(_14140_));
 OAI21_X1 _23533_ (.A(_13993_),
    .B1(_14140_),
    .B2(_13909_),
    .ZN(_14141_));
 NOR2_X2 _23534_ (.A1(_14028_),
    .A2(_13880_),
    .ZN(_14142_));
 NOR2_X2 _23535_ (.A1(_13967_),
    .A2(_13922_),
    .ZN(_14143_));
 OAI21_X1 _23536_ (.A(_14061_),
    .B1(_13923_),
    .B2(net1183),
    .ZN(_14144_));
 AOI221_X2 _23537_ (.A(_14066_),
    .B1(_14142_),
    .B2(_14143_),
    .C1(_14144_),
    .C2(_13879_),
    .ZN(_14145_));
 MUX2_X1 _23538_ (.A(_13995_),
    .B(_15024_),
    .S(_14012_),
    .Z(_14146_));
 NOR2_X2 _23539_ (.A1(_13956_),
    .A2(_13877_),
    .ZN(_14147_));
 AOI22_X1 _23540_ (.A1(_15043_),
    .A2(_14142_),
    .B1(_14120_),
    .B2(_14147_),
    .ZN(_14148_));
 OAI221_X1 _23541_ (.A(_14145_),
    .B1(_14146_),
    .B2(_14006_),
    .C1(_14088_),
    .C2(_14148_),
    .ZN(_14149_));
 OAI21_X1 _23542_ (.A(_15018_),
    .B1(_14003_),
    .B2(_14004_),
    .ZN(_14150_));
 AOI21_X4 _23543_ (.A(_13880_),
    .B1(_13957_),
    .B2(_13958_),
    .ZN(_14151_));
 BUF_X8 _23544_ (.A(_13839_),
    .Z(_14152_));
 BUF_X16 _23545_ (.A(_14152_),
    .Z(_15019_));
 AOI22_X1 _23546_ (.A1(_13985_),
    .A2(_13984_),
    .B1(_14151_),
    .B2(net1115),
    .ZN(_14153_));
 NAND4_X1 _23547_ (.A1(_13993_),
    .A2(_14133_),
    .A3(_14150_),
    .A4(_14153_),
    .ZN(_14154_));
 AND3_X1 _23548_ (.A1(_14141_),
    .A2(_14149_),
    .A3(_14154_),
    .ZN(_14155_));
 OAI21_X4 _23549_ (.A(_13985_),
    .B1(_13970_),
    .B2(_13971_),
    .ZN(_14156_));
 OAI21_X4 _23550_ (.A(_14156_),
    .B1(_14036_),
    .B2(_14046_),
    .ZN(_14157_));
 NOR2_X1 _23551_ (.A1(_13879_),
    .A2(_13924_),
    .ZN(_14158_));
 AOI21_X1 _23552_ (.A(_13898_),
    .B1(_14157_),
    .B2(_14158_),
    .ZN(_14159_));
 NAND2_X1 _23553_ (.A1(_15027_),
    .A2(_14021_),
    .ZN(_14160_));
 OAI21_X1 _23554_ (.A(_15019_),
    .B1(_14089_),
    .B2(_14003_),
    .ZN(_14161_));
 AND2_X1 _23555_ (.A1(_14160_),
    .A2(_14161_),
    .ZN(_14162_));
 AOI21_X1 _23556_ (.A(_13981_),
    .B1(_14051_),
    .B2(net1115),
    .ZN(_14163_));
 NOR2_X1 _23557_ (.A1(_14151_),
    .A2(_14163_),
    .ZN(_14164_));
 OAI221_X1 _23558_ (.A(_14159_),
    .B1(_14162_),
    .B2(_14088_),
    .C1(_15036_),
    .C2(_14164_),
    .ZN(_14165_));
 BUF_X4 _23559_ (.A(_13896_),
    .Z(_14166_));
 NAND2_X1 _23560_ (.A1(_13923_),
    .A2(_14166_),
    .ZN(_14167_));
 NOR2_X1 _23561_ (.A1(_14119_),
    .A2(_14038_),
    .ZN(_14168_));
 AOI221_X2 _23562_ (.A(_14167_),
    .B1(_14157_),
    .B2(_14119_),
    .C1(_14168_),
    .C2(_14068_),
    .ZN(_14169_));
 OAI22_X1 _23563_ (.A1(_13956_),
    .A2(_13960_),
    .B1(_14005_),
    .B2(net1115),
    .ZN(_14170_));
 NOR2_X1 _23564_ (.A1(_13924_),
    .A2(_14065_),
    .ZN(_14171_));
 AOI21_X1 _23565_ (.A(_14169_),
    .B1(_14170_),
    .B2(_14171_),
    .ZN(_14172_));
 AOI21_X1 _23566_ (.A(_14010_),
    .B1(_14165_),
    .B2(_14172_),
    .ZN(_14173_));
 OAI21_X2 _23567_ (.A(_14135_),
    .B1(_14155_),
    .B2(_14173_),
    .ZN(_00089_));
 CLKBUF_X3 _23568_ (.A(_13924_),
    .Z(_14174_));
 NAND4_X1 _23569_ (.A1(_13883_),
    .A2(_14039_),
    .A3(_14065_),
    .A4(_13968_),
    .ZN(_14175_));
 NOR2_X4 _23570_ (.A1(_14024_),
    .A2(net967),
    .ZN(_14176_));
 OR2_X1 _23571_ (.A1(_14006_),
    .A2(_14176_),
    .ZN(_14177_));
 OAI21_X1 _23572_ (.A(_14175_),
    .B1(_14177_),
    .B2(_13897_),
    .ZN(_00629_));
 CLKBUF_X3 _23573_ (.A(_14036_),
    .Z(_00630_));
 NOR2_X2 _23574_ (.A1(_13882_),
    .A2(_14166_),
    .ZN(_00631_));
 NAND2_X1 _23575_ (.A1(_00630_),
    .A2(_00631_),
    .ZN(_00632_));
 NAND2_X1 _23576_ (.A1(_13951_),
    .A2(_00631_),
    .ZN(_00633_));
 OAI22_X1 _23577_ (.A1(_14142_),
    .A2(_00632_),
    .B1(_00633_),
    .B2(_14001_),
    .ZN(_00634_));
 OAI21_X1 _23578_ (.A(_14166_),
    .B1(_14015_),
    .B2(_15048_),
    .ZN(_00635_));
 AOI21_X1 _23579_ (.A(_00635_),
    .B1(_14160_),
    .B2(_14093_),
    .ZN(_00636_));
 NOR4_X1 _23580_ (.A1(_14174_),
    .A2(_00629_),
    .A3(_00634_),
    .A4(_00636_),
    .ZN(_00637_));
 NAND2_X1 _23581_ (.A1(_13956_),
    .A2(_14003_),
    .ZN(_00638_));
 OAI21_X1 _23582_ (.A(_13883_),
    .B1(_14111_),
    .B2(_14127_),
    .ZN(_00639_));
 AOI21_X1 _23583_ (.A(_14034_),
    .B1(_00638_),
    .B2(_00639_),
    .ZN(_00640_));
 AND2_X1 _23584_ (.A1(_15039_),
    .A2(_14015_),
    .ZN(_00641_));
 NOR3_X1 _23585_ (.A1(_14029_),
    .A2(_14061_),
    .A3(_14013_),
    .ZN(_00642_));
 NOR3_X1 _23586_ (.A1(_13991_),
    .A2(_00641_),
    .A3(_00642_),
    .ZN(_00643_));
 NOR3_X1 _23587_ (.A1(_14088_),
    .A2(_00640_),
    .A3(_00643_),
    .ZN(_00644_));
 AOI21_X1 _23588_ (.A(_13998_),
    .B1(_14095_),
    .B2(_14014_),
    .ZN(_00645_));
 MUX2_X1 _23589_ (.A(_15041_),
    .B(_00645_),
    .S(_00630_),
    .Z(_00646_));
 OAI21_X1 _23590_ (.A(_13994_),
    .B1(_14129_),
    .B2(_00646_),
    .ZN(_00647_));
 NOR2_X1 _23591_ (.A1(_14028_),
    .A2(_13878_),
    .ZN(_00648_));
 NOR2_X1 _23592_ (.A1(_15024_),
    .A2(_15027_),
    .ZN(_00649_));
 NOR3_X1 _23593_ (.A1(_14108_),
    .A2(_00648_),
    .A3(_00649_),
    .ZN(_00650_));
 OAI21_X1 _23594_ (.A(_14133_),
    .B1(_14098_),
    .B2(_15044_),
    .ZN(_00651_));
 NOR2_X1 _23595_ (.A1(_00650_),
    .A2(_00651_),
    .ZN(_00652_));
 OAI21_X2 _23596_ (.A(_15028_),
    .B1(_13970_),
    .B2(_13971_),
    .ZN(_00653_));
 OAI21_X1 _23597_ (.A(_00653_),
    .B1(_14015_),
    .B2(_14014_),
    .ZN(_00654_));
 NOR3_X2 _23598_ (.A1(_13980_),
    .A2(_13945_),
    .A3(_13948_),
    .ZN(_00655_));
 OR2_X1 _23599_ (.A1(_14047_),
    .A2(_00655_),
    .ZN(_00656_));
 OAI221_X1 _23600_ (.A(_14171_),
    .B1(_00654_),
    .B2(_13879_),
    .C1(_00656_),
    .C2(net1188),
    .ZN(_00657_));
 MUX2_X1 _23601_ (.A(_14020_),
    .B(_13950_),
    .S(_13840_),
    .Z(_00658_));
 AOI222_X2 _23602_ (.A1(_14042_),
    .A2(_14059_),
    .B1(_13976_),
    .B2(_00648_),
    .C1(_00658_),
    .C2(_13985_),
    .ZN(_00659_));
 NAND2_X2 _23603_ (.A1(_14012_),
    .A2(_13991_),
    .ZN(_00660_));
 OAI21_X1 _23604_ (.A(_00657_),
    .B1(_00659_),
    .B2(_00660_),
    .ZN(_00661_));
 OAI33_X1 _23605_ (.A1(_14010_),
    .A2(_00637_),
    .A3(_00644_),
    .B1(_00647_),
    .B2(_00652_),
    .B3(_00661_),
    .ZN(_00662_));
 OR4_X1 _23606_ (.A1(_14028_),
    .A2(_13881_),
    .A3(_14078_),
    .A4(_14073_),
    .ZN(_00663_));
 AOI21_X1 _23607_ (.A(_14011_),
    .B1(_14113_),
    .B2(_14117_),
    .ZN(_00664_));
 OAI21_X1 _23608_ (.A(_14047_),
    .B1(_13996_),
    .B2(_14151_),
    .ZN(_00665_));
 OAI21_X1 _23609_ (.A(_13878_),
    .B1(_14018_),
    .B2(_14024_),
    .ZN(_00666_));
 NOR2_X1 _23610_ (.A1(net960),
    .A2(_14036_),
    .ZN(_00667_));
 OAI21_X1 _23611_ (.A(_00665_),
    .B1(_00666_),
    .B2(_00667_),
    .ZN(_00668_));
 AOI221_X2 _23612_ (.A(_13897_),
    .B1(_00663_),
    .B2(_00664_),
    .C1(_00668_),
    .C2(_14012_),
    .ZN(_00669_));
 OAI22_X2 _23613_ (.A1(_13956_),
    .A2(_13882_),
    .B1(_14099_),
    .B2(_14028_),
    .ZN(_00670_));
 AOI221_X2 _23614_ (.A(_14011_),
    .B1(_14057_),
    .B2(_14058_),
    .C1(_00670_),
    .C2(_14015_),
    .ZN(_00671_));
 MUX2_X1 _23615_ (.A(_14017_),
    .B(_15025_),
    .S(_13881_),
    .Z(_00672_));
 OAI21_X2 _23616_ (.A(_13964_),
    .B1(_14061_),
    .B2(_00672_),
    .ZN(_00673_));
 AOI21_X2 _23617_ (.A(_00673_),
    .B1(_14160_),
    .B2(_14093_),
    .ZN(_00674_));
 NOR3_X2 _23618_ (.A1(_00671_),
    .A2(_00674_),
    .A3(_13992_),
    .ZN(_00675_));
 NOR3_X4 _23619_ (.A1(_14117_),
    .A2(_13970_),
    .A3(_13971_),
    .ZN(_00676_));
 NOR2_X2 _23620_ (.A1(_14137_),
    .A2(_00676_),
    .ZN(_00677_));
 OAI221_X2 _23621_ (.A(_14011_),
    .B1(_14059_),
    .B2(_13950_),
    .C1(_00677_),
    .C2(_13882_),
    .ZN(_00678_));
 NAND2_X1 _23622_ (.A1(_13956_),
    .A2(_13965_),
    .ZN(_00679_));
 NAND3_X1 _23623_ (.A1(_13840_),
    .A2(_13881_),
    .A3(_13967_),
    .ZN(_00680_));
 NAND3_X1 _23624_ (.A1(_13923_),
    .A2(_00679_),
    .A3(_00680_),
    .ZN(_00681_));
 AOI221_X2 _23625_ (.A(_14065_),
    .B1(_00678_),
    .B2(_00681_),
    .C1(_14004_),
    .C2(_13952_),
    .ZN(_00682_));
 NOR2_X4 _23626_ (.A1(_13877_),
    .A2(_13941_),
    .ZN(_00683_));
 OAI21_X1 _23627_ (.A(_14120_),
    .B1(_14015_),
    .B2(_13953_),
    .ZN(_00684_));
 AOI221_X2 _23628_ (.A(_14129_),
    .B1(_00683_),
    .B2(_13981_),
    .C1(_00684_),
    .C2(_14119_),
    .ZN(_00685_));
 AOI21_X1 _23629_ (.A(_14089_),
    .B1(_14061_),
    .B2(_13952_),
    .ZN(_00686_));
 NOR2_X1 _23630_ (.A1(_13883_),
    .A2(_00676_),
    .ZN(_00687_));
 NAND2_X1 _23631_ (.A1(_14152_),
    .A2(_14061_),
    .ZN(_00688_));
 AOI22_X1 _23632_ (.A1(_13883_),
    .A2(_00686_),
    .B1(_00687_),
    .B2(_00688_),
    .ZN(_00689_));
 OAI21_X1 _23633_ (.A(_13994_),
    .B1(_00660_),
    .B2(_00689_),
    .ZN(_00690_));
 OAI33_X1 _23634_ (.A1(_00675_),
    .A2(_00669_),
    .A3(_14010_),
    .B1(_00682_),
    .B2(_00685_),
    .B3(_00690_),
    .ZN(_00691_));
 MUX2_X1 _23635_ (.A(_00662_),
    .B(_00691_),
    .S(_14104_),
    .Z(_00090_));
 NOR2_X1 _23636_ (.A1(_14010_),
    .A2(_13898_),
    .ZN(_00692_));
 NAND2_X1 _23637_ (.A1(_14001_),
    .A2(_14039_),
    .ZN(_00693_));
 AOI21_X1 _23638_ (.A(_13879_),
    .B1(_00630_),
    .B2(net572),
    .ZN(_00694_));
 NAND2_X1 _23639_ (.A1(_00693_),
    .A2(_00694_),
    .ZN(_00695_));
 OAI21_X1 _23640_ (.A(_15043_),
    .B1(_14089_),
    .B2(_13941_),
    .ZN(_00696_));
 NAND4_X1 _23641_ (.A1(_14088_),
    .A2(_13993_),
    .A3(_00695_),
    .A4(_00696_),
    .ZN(_00697_));
 NOR3_X1 _23642_ (.A1(_15043_),
    .A2(_14038_),
    .A3(net1206),
    .ZN(_00698_));
 AOI21_X1 _23643_ (.A(_14054_),
    .B1(_14108_),
    .B2(net1115),
    .ZN(_00699_));
 AOI21_X1 _23644_ (.A(_00698_),
    .B1(_00699_),
    .B2(_15043_),
    .ZN(_00700_));
 NAND3_X1 _23645_ (.A1(_14174_),
    .A2(_13993_),
    .A3(_00700_),
    .ZN(_00701_));
 NAND2_X1 _23646_ (.A1(_13883_),
    .A2(_13964_),
    .ZN(_00702_));
 AOI21_X1 _23647_ (.A(_14081_),
    .B1(_14098_),
    .B2(_14024_),
    .ZN(_00703_));
 AOI22_X1 _23648_ (.A1(_14108_),
    .A2(_14026_),
    .B1(_14005_),
    .B2(_13952_),
    .ZN(_00704_));
 OAI221_X1 _23649_ (.A(_14104_),
    .B1(_00702_),
    .B2(_00703_),
    .C1(_00704_),
    .C2(_14088_),
    .ZN(_00705_));
 NAND4_X1 _23650_ (.A1(_00692_),
    .A2(_00697_),
    .A3(_00701_),
    .A4(_00705_),
    .ZN(_00706_));
 NAND2_X1 _23651_ (.A1(_13909_),
    .A2(_13898_),
    .ZN(_00707_));
 AOI21_X1 _23652_ (.A(_14104_),
    .B1(_14158_),
    .B2(_15027_),
    .ZN(_00708_));
 NOR3_X1 _23653_ (.A1(net1115),
    .A2(_15036_),
    .A3(_14043_),
    .ZN(_00709_));
 NOR3_X1 _23654_ (.A1(net1187),
    .A2(_14012_),
    .A3(_14026_),
    .ZN(_00710_));
 NOR3_X1 _23655_ (.A1(_14098_),
    .A2(_00709_),
    .A3(_00710_),
    .ZN(_00711_));
 NOR3_X1 _23656_ (.A1(_14029_),
    .A2(_13883_),
    .A3(_13964_),
    .ZN(_00712_));
 AOI21_X1 _23657_ (.A(_13995_),
    .B1(_13879_),
    .B2(_13924_),
    .ZN(_00713_));
 NOR4_X1 _23658_ (.A1(_14108_),
    .A2(_14158_),
    .A3(_00712_),
    .A4(_00713_),
    .ZN(_00714_));
 OAI21_X1 _23659_ (.A(_00708_),
    .B1(_00711_),
    .B2(_00714_),
    .ZN(_00715_));
 NAND2_X1 _23660_ (.A1(net1185),
    .A2(_14018_),
    .ZN(_00716_));
 AOI21_X1 _23661_ (.A(_14111_),
    .B1(_13951_),
    .B2(_14001_),
    .ZN(_00717_));
 AOI221_X2 _23662_ (.A(_13924_),
    .B1(_00716_),
    .B2(_14070_),
    .C1(_00717_),
    .C2(_14119_),
    .ZN(_00718_));
 NOR3_X2 _23663_ (.A1(_14047_),
    .A2(_14038_),
    .A3(_14067_),
    .ZN(_00719_));
 AOI21_X1 _23664_ (.A(_14081_),
    .B1(_14176_),
    .B2(_14098_),
    .ZN(_00720_));
 AOI21_X1 _23665_ (.A(_00719_),
    .B1(_00720_),
    .B2(_15036_),
    .ZN(_00721_));
 AOI21_X1 _23666_ (.A(_00718_),
    .B1(_00721_),
    .B2(_14174_),
    .ZN(_00722_));
 OAI21_X1 _23667_ (.A(_00715_),
    .B1(_00722_),
    .B2(_13993_),
    .ZN(_00723_));
 MUX2_X1 _23668_ (.A(_13953_),
    .B(_14176_),
    .S(_14047_),
    .Z(_00724_));
 OAI21_X1 _23669_ (.A(_14107_),
    .B1(_00724_),
    .B2(_14108_),
    .ZN(_00725_));
 AOI21_X1 _23670_ (.A(_14026_),
    .B1(_14119_),
    .B2(net1183),
    .ZN(_00726_));
 AOI21_X1 _23671_ (.A(_13991_),
    .B1(_14143_),
    .B2(_00726_),
    .ZN(_00727_));
 AOI21_X1 _23672_ (.A(_13965_),
    .B1(_14018_),
    .B2(_14028_),
    .ZN(_00728_));
 OAI221_X2 _23673_ (.A(_14114_),
    .B1(_00728_),
    .B2(_15018_),
    .C1(_13960_),
    .C2(_14029_),
    .ZN(_00729_));
 AOI21_X4 _23674_ (.A(_15030_),
    .B1(_13957_),
    .B2(_13958_),
    .ZN(_00730_));
 NOR2_X1 _23675_ (.A1(_14081_),
    .A2(_00730_),
    .ZN(_00731_));
 NOR3_X4 _23676_ (.A1(_14017_),
    .A2(_13970_),
    .A3(_13971_),
    .ZN(_00732_));
 NOR2_X1 _23677_ (.A1(_14151_),
    .A2(_00732_),
    .ZN(_00733_));
 MUX2_X1 _23678_ (.A(_00731_),
    .B(_00733_),
    .S(_13878_),
    .Z(_00734_));
 MUX2_X1 _23679_ (.A(_00729_),
    .B(_00734_),
    .S(_14012_),
    .Z(_00735_));
 AOI221_X2 _23680_ (.A(_13993_),
    .B1(_00725_),
    .B2(_00727_),
    .C1(_00735_),
    .C2(_13992_),
    .ZN(_00736_));
 AOI221_X1 _23681_ (.A(_14129_),
    .B1(_14113_),
    .B2(_14001_),
    .C1(_13995_),
    .C2(_13984_),
    .ZN(_00737_));
 AOI22_X1 _23682_ (.A1(_14108_),
    .A2(_14026_),
    .B1(_14003_),
    .B2(_15018_),
    .ZN(_00738_));
 OAI21_X1 _23683_ (.A(_00737_),
    .B1(_00738_),
    .B2(net1115),
    .ZN(_00739_));
 NAND2_X2 _23684_ (.A1(_14028_),
    .A2(_14073_),
    .ZN(_00740_));
 NAND3_X1 _23685_ (.A1(_14002_),
    .A2(_00665_),
    .A3(_00740_),
    .ZN(_00741_));
 OAI21_X1 _23686_ (.A(_00739_),
    .B1(_00741_),
    .B2(_00660_),
    .ZN(_00742_));
 AOI211_X2 _23687_ (.A(_14020_),
    .B(_13996_),
    .C1(_14036_),
    .C2(_14028_),
    .ZN(_00743_));
 AOI21_X1 _23688_ (.A(_14038_),
    .B1(_14039_),
    .B2(_13953_),
    .ZN(_00744_));
 AOI21_X1 _23689_ (.A(_00743_),
    .B1(_00744_),
    .B2(_15043_),
    .ZN(_00745_));
 NOR3_X1 _23690_ (.A1(_14113_),
    .A2(_00649_),
    .A3(_14094_),
    .ZN(_00746_));
 OAI221_X1 _23691_ (.A(_13993_),
    .B1(_14136_),
    .B2(_00745_),
    .C1(_00746_),
    .C2(_14167_),
    .ZN(_00747_));
 OAI21_X1 _23692_ (.A(_14010_),
    .B1(_00747_),
    .B2(_00742_),
    .ZN(_00748_));
 OAI221_X1 _23693_ (.A(_00706_),
    .B1(_00707_),
    .B2(_00723_),
    .C1(_00736_),
    .C2(_00748_),
    .ZN(_00091_));
 NAND2_X1 _23694_ (.A1(_13994_),
    .A2(_13902_),
    .ZN(_00749_));
 AOI21_X1 _23695_ (.A(_13883_),
    .B1(_00630_),
    .B2(_13952_),
    .ZN(_00750_));
 OAI21_X1 _23696_ (.A(_14031_),
    .B1(_14053_),
    .B2(_00750_),
    .ZN(_00751_));
 OAI221_X1 _23697_ (.A(_14051_),
    .B1(_14093_),
    .B2(_00656_),
    .C1(_14022_),
    .C2(_15018_),
    .ZN(_00752_));
 AND3_X1 _23698_ (.A1(_13992_),
    .A2(_00751_),
    .A3(_00752_),
    .ZN(_00753_));
 AOI21_X1 _23699_ (.A(_13859_),
    .B1(_13965_),
    .B2(_13922_),
    .ZN(_00754_));
 OAI221_X2 _23700_ (.A(_13951_),
    .B1(_00754_),
    .B2(net960),
    .C1(_15018_),
    .C2(_14021_),
    .ZN(_00755_));
 MUX2_X1 _23701_ (.A(_14057_),
    .B(_14100_),
    .S(_13963_),
    .Z(_00756_));
 NAND2_X1 _23702_ (.A1(_00630_),
    .A2(_00756_),
    .ZN(_00757_));
 OAI21_X1 _23703_ (.A(_00702_),
    .B1(_14045_),
    .B2(_15027_),
    .ZN(_00758_));
 AOI221_X2 _23704_ (.A(_13991_),
    .B1(_00755_),
    .B2(_00757_),
    .C1(_00758_),
    .C2(net1115),
    .ZN(_00759_));
 NOR3_X1 _23705_ (.A1(_00749_),
    .A2(_00753_),
    .A3(_00759_),
    .ZN(_00760_));
 NOR3_X1 _23706_ (.A1(net967),
    .A2(_13970_),
    .A3(_13971_),
    .ZN(_00761_));
 NOR2_X2 _23707_ (.A1(_13965_),
    .A2(_00761_),
    .ZN(_00762_));
 OAI21_X1 _23708_ (.A(_00762_),
    .B1(_13976_),
    .B2(_14152_),
    .ZN(_00763_));
 NOR3_X1 _23709_ (.A1(_13882_),
    .A2(_14073_),
    .A3(_13996_),
    .ZN(_00764_));
 NOR2_X1 _23710_ (.A1(_14166_),
    .A2(_00764_),
    .ZN(_00765_));
 OAI22_X1 _23711_ (.A1(net1183),
    .A2(_13960_),
    .B1(_14067_),
    .B2(_14119_),
    .ZN(_00766_));
 AOI221_X2 _23712_ (.A(_14012_),
    .B1(_00763_),
    .B2(_00765_),
    .C1(_00766_),
    .C2(_14034_),
    .ZN(_00767_));
 NOR3_X1 _23713_ (.A1(_14020_),
    .A2(_14054_),
    .A3(_00655_),
    .ZN(_00768_));
 AOI21_X1 _23714_ (.A(_00768_),
    .B1(_14091_),
    .B2(_14021_),
    .ZN(_00769_));
 OAI22_X1 _23715_ (.A1(_14024_),
    .A2(_14061_),
    .B1(_13976_),
    .B2(net960),
    .ZN(_00770_));
 AOI221_X2 _23716_ (.A(_14051_),
    .B1(_13897_),
    .B2(_00769_),
    .C1(_00770_),
    .C2(_00631_),
    .ZN(_00771_));
 NOR3_X2 _23717_ (.A1(_14126_),
    .A2(_00767_),
    .A3(_00771_),
    .ZN(_00772_));
 NAND2_X1 _23718_ (.A1(_13909_),
    .A2(_13902_),
    .ZN(_00773_));
 NOR2_X1 _23719_ (.A1(_14021_),
    .A2(_00732_),
    .ZN(_00774_));
 AOI221_X1 _23720_ (.A(_14129_),
    .B1(_00731_),
    .B2(_14021_),
    .C1(_00774_),
    .C2(_14074_),
    .ZN(_00775_));
 MUX2_X1 _23721_ (.A(_13956_),
    .B(_14014_),
    .S(_14015_),
    .Z(_00776_));
 AOI22_X1 _23722_ (.A1(_14068_),
    .A2(_00694_),
    .B1(_00776_),
    .B2(_14022_),
    .ZN(_00777_));
 AOI21_X1 _23723_ (.A(_00775_),
    .B1(_00777_),
    .B2(_14133_),
    .ZN(_00778_));
 AOI21_X2 _23724_ (.A(_00732_),
    .B1(_14036_),
    .B2(net960),
    .ZN(_00779_));
 AOI22_X2 _23725_ (.A1(_14074_),
    .A2(_00762_),
    .B1(_00779_),
    .B2(_14022_),
    .ZN(_00780_));
 OAI21_X1 _23726_ (.A(_13991_),
    .B1(_15043_),
    .B2(_13952_),
    .ZN(_00781_));
 NOR2_X1 _23727_ (.A1(_15036_),
    .A2(_14157_),
    .ZN(_00782_));
 OAI221_X2 _23728_ (.A(_14088_),
    .B1(_13992_),
    .B2(_00780_),
    .C1(_00782_),
    .C2(_00781_),
    .ZN(_00783_));
 AOI21_X2 _23729_ (.A(_00773_),
    .B1(_00783_),
    .B2(_00778_),
    .ZN(_00784_));
 NOR2_X1 _23730_ (.A1(_14061_),
    .A2(_14166_),
    .ZN(_00785_));
 OAI21_X1 _23731_ (.A(_13879_),
    .B1(_00730_),
    .B2(_00785_),
    .ZN(_00786_));
 NAND3_X1 _23732_ (.A1(_13859_),
    .A2(_14113_),
    .A3(_13896_),
    .ZN(_00787_));
 NAND3_X1 _23733_ (.A1(_14011_),
    .A2(_14068_),
    .A3(_00787_),
    .ZN(_00788_));
 OAI21_X1 _23734_ (.A(_13960_),
    .B1(_14166_),
    .B2(_14006_),
    .ZN(_00789_));
 AOI21_X1 _23735_ (.A(_00788_),
    .B1(_00789_),
    .B2(_14029_),
    .ZN(_00790_));
 OAI221_X1 _23736_ (.A(_00740_),
    .B1(_13977_),
    .B2(_13965_),
    .C1(_15020_),
    .C2(_13960_),
    .ZN(_00791_));
 OAI21_X1 _23737_ (.A(_13967_),
    .B1(_13882_),
    .B2(_13995_),
    .ZN(_00792_));
 OAI21_X1 _23738_ (.A(_00792_),
    .B1(_14015_),
    .B2(_15032_),
    .ZN(_00793_));
 MUX2_X1 _23739_ (.A(_00791_),
    .B(_00793_),
    .S(_14065_),
    .Z(_00794_));
 AOI221_X2 _23740_ (.A(_14105_),
    .B1(_00786_),
    .B2(_00790_),
    .C1(_00794_),
    .C2(_14051_),
    .ZN(_00795_));
 NOR4_X2 _23741_ (.A1(_00784_),
    .A2(_00772_),
    .A3(_00760_),
    .A4(_00795_),
    .ZN(_00092_));
 OAI221_X1 _23742_ (.A(_13897_),
    .B1(_13969_),
    .B2(_13973_),
    .C1(_14059_),
    .C2(_00630_),
    .ZN(_00796_));
 OAI221_X1 _23743_ (.A(_14065_),
    .B1(_13981_),
    .B2(_14029_),
    .C1(_14004_),
    .C2(_15018_),
    .ZN(_00797_));
 AND3_X1 _23744_ (.A1(_14051_),
    .A2(_00796_),
    .A3(_00797_),
    .ZN(_00798_));
 OAI21_X1 _23745_ (.A(_14121_),
    .B1(_13950_),
    .B2(_14001_),
    .ZN(_00799_));
 AOI22_X2 _23746_ (.A1(_13968_),
    .A2(_14004_),
    .B1(_00799_),
    .B2(_14022_),
    .ZN(_00800_));
 AOI21_X1 _23747_ (.A(_14047_),
    .B1(_13951_),
    .B2(_13953_),
    .ZN(_00801_));
 AOI22_X2 _23748_ (.A1(_13999_),
    .A2(_00683_),
    .B1(_00801_),
    .B2(_14074_),
    .ZN(_00802_));
 OAI22_X2 _23749_ (.A1(_14136_),
    .A2(_00800_),
    .B1(_00802_),
    .B2(_00660_),
    .ZN(_00803_));
 OR3_X2 _23750_ (.A1(_14126_),
    .A2(_00798_),
    .A3(_00803_),
    .ZN(_00804_));
 OAI221_X1 _23751_ (.A(_14031_),
    .B1(_13972_),
    .B2(_14071_),
    .C1(_14099_),
    .C2(_14098_),
    .ZN(_00805_));
 OAI21_X1 _23752_ (.A(_14051_),
    .B1(_13984_),
    .B2(net1187),
    .ZN(_00806_));
 AOI21_X1 _23753_ (.A(_13898_),
    .B1(_00805_),
    .B2(_00806_),
    .ZN(_00807_));
 OAI21_X1 _23754_ (.A(_15027_),
    .B1(_14143_),
    .B2(net1187),
    .ZN(_00808_));
 OAI21_X1 _23755_ (.A(net1187),
    .B1(_00630_),
    .B2(_14012_),
    .ZN(_00809_));
 AOI21_X1 _23756_ (.A(_00809_),
    .B1(_14113_),
    .B2(_14031_),
    .ZN(_00810_));
 OAI21_X1 _23757_ (.A(_00807_),
    .B1(_00808_),
    .B2(_00810_),
    .ZN(_00811_));
 AND2_X2 _23758_ (.A1(_13975_),
    .A2(_14156_),
    .ZN(_00812_));
 OAI221_X1 _23759_ (.A(_14031_),
    .B1(_14025_),
    .B2(net1187),
    .C1(_00812_),
    .C2(_15036_),
    .ZN(_00813_));
 AOI21_X1 _23760_ (.A(_00676_),
    .B1(_14098_),
    .B2(_13980_),
    .ZN(_00814_));
 OAI221_X1 _23761_ (.A(_14174_),
    .B1(_14006_),
    .B2(_13985_),
    .C1(_00814_),
    .C2(_15036_),
    .ZN(_00815_));
 NAND3_X1 _23762_ (.A1(_00813_),
    .A2(_13898_),
    .A3(_00815_),
    .ZN(_00816_));
 NAND4_X2 _23763_ (.A1(_00816_),
    .A2(_13993_),
    .A3(_00811_),
    .A4(_13909_),
    .ZN(_00817_));
 AOI22_X2 _23764_ (.A1(_13956_),
    .A2(_13950_),
    .B1(_14074_),
    .B2(_14020_),
    .ZN(_00818_));
 NAND2_X1 _23765_ (.A1(_15030_),
    .A2(_13876_),
    .ZN(_00819_));
 NOR2_X1 _23766_ (.A1(_13967_),
    .A2(_00819_),
    .ZN(_00820_));
 NOR3_X1 _23767_ (.A1(_14166_),
    .A2(_14137_),
    .A3(_00820_),
    .ZN(_00821_));
 NAND2_X1 _23768_ (.A1(_14068_),
    .A2(_14070_),
    .ZN(_00822_));
 AOI221_X2 _23769_ (.A(_13924_),
    .B1(_14166_),
    .B2(_00818_),
    .C1(_00821_),
    .C2(_00822_),
    .ZN(_00823_));
 OAI221_X1 _23770_ (.A(_14133_),
    .B1(_00731_),
    .B2(_13879_),
    .C1(_13972_),
    .C2(_15018_),
    .ZN(_00824_));
 AND2_X4 _23771_ (.A1(_00672_),
    .A2(_14015_),
    .ZN(_00825_));
 MUX2_X1 _23772_ (.A(_14024_),
    .B(net960),
    .S(_13878_),
    .Z(_00826_));
 AOI21_X4 _23773_ (.A(_00825_),
    .B1(_00826_),
    .B2(_14108_),
    .ZN(_00827_));
 OAI21_X4 _23774_ (.A(_00824_),
    .B1(_00827_),
    .B2(_14129_),
    .ZN(_00828_));
 OR3_X4 _23775_ (.A1(_00828_),
    .A2(_00823_),
    .A3(_00749_),
    .ZN(_00829_));
 NAND2_X2 _23776_ (.A1(_13985_),
    .A2(_13950_),
    .ZN(_00830_));
 AOI221_X2 _23777_ (.A(_13990_),
    .B1(_00683_),
    .B2(_00830_),
    .C1(_00799_),
    .C2(_13878_),
    .ZN(_00831_));
 NAND2_X1 _23778_ (.A1(_14117_),
    .A2(_13965_),
    .ZN(_00832_));
 AOI221_X1 _23779_ (.A(_14166_),
    .B1(_13984_),
    .B2(_13956_),
    .C1(_00832_),
    .C2(_14036_),
    .ZN(_00833_));
 OR3_X2 _23780_ (.A1(_00831_),
    .A2(_14174_),
    .A3(_00833_),
    .ZN(_00834_));
 AOI221_X2 _23781_ (.A(_13897_),
    .B1(_14176_),
    .B2(_14113_),
    .C1(_14096_),
    .C2(_00667_),
    .ZN(_00835_));
 AOI221_X1 _23782_ (.A(_14065_),
    .B1(_14142_),
    .B2(_14004_),
    .C1(_00630_),
    .C2(_14001_),
    .ZN(_00836_));
 OAI21_X1 _23783_ (.A(_14174_),
    .B1(_00835_),
    .B2(_00836_),
    .ZN(_00837_));
 NAND4_X4 _23784_ (.A1(_13909_),
    .A2(_14104_),
    .A3(_00834_),
    .A4(_00837_),
    .ZN(_00838_));
 AND4_X4 _23785_ (.A1(_00838_),
    .A2(_00817_),
    .A3(_00804_),
    .A4(_00829_),
    .ZN(_00093_));
 NAND2_X1 _23786_ (.A1(_13953_),
    .A2(_14036_),
    .ZN(_00839_));
 NOR2_X1 _23787_ (.A1(_13877_),
    .A2(_00655_),
    .ZN(_00840_));
 AOI221_X2 _23788_ (.A(_13897_),
    .B1(_00839_),
    .B2(_00840_),
    .C1(_14003_),
    .C2(_14024_),
    .ZN(_00841_));
 NOR3_X1 _23789_ (.A1(_14022_),
    .A2(_14089_),
    .A3(_00730_),
    .ZN(_00842_));
 AOI21_X1 _23790_ (.A(net1206),
    .B1(_14176_),
    .B2(_14098_),
    .ZN(_00843_));
 AOI21_X1 _23791_ (.A(_00842_),
    .B1(_00843_),
    .B2(_15043_),
    .ZN(_00844_));
 AOI21_X1 _23792_ (.A(_00841_),
    .B1(_00844_),
    .B2(_13898_),
    .ZN(_00845_));
 NOR3_X1 _23793_ (.A1(_00845_),
    .A2(_14174_),
    .A3(_13909_),
    .ZN(_00846_));
 AOI21_X1 _23794_ (.A(_14021_),
    .B1(_14061_),
    .B2(_14024_),
    .ZN(_00847_));
 OAI22_X1 _23795_ (.A1(_13952_),
    .A2(_00630_),
    .B1(_13976_),
    .B2(_14029_),
    .ZN(_00848_));
 AOI221_X2 _23796_ (.A(_13991_),
    .B1(_14121_),
    .B2(_00847_),
    .C1(_00848_),
    .C2(_14022_),
    .ZN(_00849_));
 OAI221_X2 _23797_ (.A(_13968_),
    .B1(_13971_),
    .B2(_13970_),
    .C1(net1185),
    .C2(_14020_),
    .ZN(_00850_));
 OR3_X1 _23798_ (.A1(_15037_),
    .A2(_15046_),
    .A3(_00630_),
    .ZN(_00851_));
 NAND3_X1 _23799_ (.A1(_13992_),
    .A2(_00850_),
    .A3(_00851_),
    .ZN(_00852_));
 NAND3_X1 _23800_ (.A1(_14010_),
    .A2(_14174_),
    .A3(_00852_),
    .ZN(_00853_));
 OAI21_X1 _23801_ (.A(_13993_),
    .B1(_00849_),
    .B2(_00853_),
    .ZN(_00854_));
 OR2_X1 _23802_ (.A1(_15039_),
    .A2(_13951_),
    .ZN(_00855_));
 OAI221_X1 _23803_ (.A(_14039_),
    .B1(_14013_),
    .B2(_14152_),
    .C1(_14119_),
    .C2(_13985_),
    .ZN(_00856_));
 NAND3_X1 _23804_ (.A1(_13991_),
    .A2(_00855_),
    .A3(_00856_),
    .ZN(_00857_));
 NOR2_X1 _23805_ (.A1(_14029_),
    .A2(_14026_),
    .ZN(_00858_));
 OAI221_X1 _23806_ (.A(_14034_),
    .B1(_13960_),
    .B2(_14001_),
    .C1(_00858_),
    .C2(_14108_),
    .ZN(_00859_));
 AND3_X1 _23807_ (.A1(_14031_),
    .A2(_00857_),
    .A3(_00859_),
    .ZN(_00860_));
 AOI21_X1 _23808_ (.A(_14020_),
    .B1(_13950_),
    .B2(_14176_),
    .ZN(_00861_));
 NOR2_X1 _23809_ (.A1(_13996_),
    .A2(_14151_),
    .ZN(_00862_));
 AOI221_X1 _23810_ (.A(_14065_),
    .B1(_14074_),
    .B2(_00861_),
    .C1(_00862_),
    .C2(_14021_),
    .ZN(_00863_));
 AOI221_X2 _23811_ (.A(_13882_),
    .B1(_13950_),
    .B2(_14069_),
    .C1(_14073_),
    .C2(net1185),
    .ZN(_00864_));
 NOR3_X1 _23812_ (.A1(_00743_),
    .A2(_14034_),
    .A3(_00864_),
    .ZN(_00865_));
 NOR3_X1 _23813_ (.A1(_00865_),
    .A2(_00863_),
    .A3(_14088_),
    .ZN(_00866_));
 NOR3_X1 _23814_ (.A1(_14010_),
    .A2(_00860_),
    .A3(_00866_),
    .ZN(_00867_));
 NAND2_X1 _23815_ (.A1(_13994_),
    .A2(_14166_),
    .ZN(_00868_));
 MUX2_X1 _23816_ (.A(_14028_),
    .B(_14073_),
    .S(_13922_),
    .Z(_00869_));
 AOI221_X2 _23817_ (.A(_00868_),
    .B1(_00869_),
    .B2(_14119_),
    .C1(_14012_),
    .C2(_14089_),
    .ZN(_00870_));
 AOI21_X1 _23818_ (.A(_14108_),
    .B1(_14051_),
    .B2(_13953_),
    .ZN(_00871_));
 AOI21_X1 _23819_ (.A(_00871_),
    .B1(net1206),
    .B2(_14174_),
    .ZN(_00872_));
 OAI21_X1 _23820_ (.A(_00870_),
    .B1(_00872_),
    .B2(_15043_),
    .ZN(_00873_));
 NAND2_X1 _23821_ (.A1(_14104_),
    .A2(_00873_),
    .ZN(_00874_));
 AOI21_X1 _23822_ (.A(_00719_),
    .B1(_14113_),
    .B2(_13995_),
    .ZN(_00875_));
 AOI21_X1 _23823_ (.A(_15036_),
    .B1(_00693_),
    .B2(_00839_),
    .ZN(_00876_));
 OAI21_X1 _23824_ (.A(_14034_),
    .B1(_14006_),
    .B2(net1187),
    .ZN(_00877_));
 OAI221_X1 _23825_ (.A(_14088_),
    .B1(_13898_),
    .B2(_00875_),
    .C1(_00876_),
    .C2(_00877_),
    .ZN(_00878_));
 NAND2_X1 _23826_ (.A1(_15038_),
    .A2(_14098_),
    .ZN(_00879_));
 NAND3_X1 _23827_ (.A1(_14039_),
    .A2(_14057_),
    .A3(_00819_),
    .ZN(_00880_));
 AOI21_X1 _23828_ (.A(_14034_),
    .B1(_00879_),
    .B2(_00880_),
    .ZN(_00881_));
 AND3_X1 _23829_ (.A1(_14098_),
    .A2(_13897_),
    .A3(_00670_),
    .ZN(_00882_));
 OAI21_X1 _23830_ (.A(_14174_),
    .B1(_00881_),
    .B2(_00882_),
    .ZN(_00883_));
 AOI21_X1 _23831_ (.A(_14010_),
    .B1(_00878_),
    .B2(_00883_),
    .ZN(_00884_));
 NOR2_X1 _23832_ (.A1(_14045_),
    .A2(_14059_),
    .ZN(_00885_));
 OAI21_X1 _23833_ (.A(_13882_),
    .B1(_13922_),
    .B2(_00732_),
    .ZN(_00886_));
 OAI21_X1 _23834_ (.A(_00886_),
    .B1(_14011_),
    .B2(_15027_),
    .ZN(_00887_));
 AOI21_X1 _23835_ (.A(_14078_),
    .B1(_14095_),
    .B2(net149),
    .ZN(_00888_));
 OAI221_X2 _23836_ (.A(_00740_),
    .B1(_00888_),
    .B2(net1183),
    .C1(_13880_),
    .C2(_14047_),
    .ZN(_00889_));
 AOI221_X2 _23837_ (.A(_00885_),
    .B1(_00887_),
    .B2(_14014_),
    .C1(_13964_),
    .C2(_00889_),
    .ZN(_00890_));
 NOR3_X1 _23838_ (.A1(_13909_),
    .A2(_13898_),
    .A3(_00890_),
    .ZN(_00891_));
 OAI33_X1 _23839_ (.A1(_00846_),
    .A2(_00867_),
    .A3(_00854_),
    .B1(_00874_),
    .B2(_00884_),
    .B3(_00891_),
    .ZN(_00094_));
 OAI221_X2 _23840_ (.A(_14065_),
    .B1(_13972_),
    .B2(_13952_),
    .C1(_00779_),
    .C2(_14119_),
    .ZN(_00892_));
 NOR2_X1 _23841_ (.A1(_13949_),
    .A2(_13990_),
    .ZN(_00893_));
 OAI21_X1 _23842_ (.A(_14059_),
    .B1(_13881_),
    .B2(net149),
    .ZN(_00894_));
 OAI21_X1 _23843_ (.A(_00819_),
    .B1(_14020_),
    .B2(_14117_),
    .ZN(_00895_));
 AOI221_X1 _23844_ (.A(_13963_),
    .B1(_00893_),
    .B2(_00894_),
    .C1(_00895_),
    .C2(_14018_),
    .ZN(_00896_));
 OAI221_X1 _23845_ (.A(_13990_),
    .B1(_13959_),
    .B2(_13859_),
    .C1(_14006_),
    .C2(_13980_),
    .ZN(_00897_));
 OAI21_X1 _23846_ (.A(_13981_),
    .B1(_13972_),
    .B2(_13880_),
    .ZN(_00898_));
 AOI21_X1 _23847_ (.A(_00897_),
    .B1(_00898_),
    .B2(net1187),
    .ZN(_00899_));
 OAI222_X2 _23848_ (.A1(_14117_),
    .A2(_14006_),
    .B1(_13960_),
    .B2(_15018_),
    .C1(_14005_),
    .C2(_13995_),
    .ZN(_00900_));
 AOI21_X1 _23849_ (.A(_00899_),
    .B1(_00900_),
    .B2(_14034_),
    .ZN(_00901_));
 AOI221_X1 _23850_ (.A(_14126_),
    .B1(_00892_),
    .B2(_00896_),
    .C1(_00901_),
    .C2(_14031_),
    .ZN(_00902_));
 AOI21_X1 _23851_ (.A(_14147_),
    .B1(_13878_),
    .B2(_14152_),
    .ZN(_00903_));
 OAI221_X2 _23852_ (.A(_13964_),
    .B1(_00716_),
    .B2(_14026_),
    .C1(_00903_),
    .C2(_13951_),
    .ZN(_00904_));
 NAND3_X1 _23853_ (.A1(_14024_),
    .A2(_14020_),
    .A3(_13950_),
    .ZN(_00905_));
 OAI21_X1 _23854_ (.A(_00905_),
    .B1(_14018_),
    .B2(_15032_),
    .ZN(_00906_));
 AOI21_X1 _23855_ (.A(_13897_),
    .B1(_00906_),
    .B2(_13923_),
    .ZN(_00907_));
 OAI21_X1 _23856_ (.A(_13923_),
    .B1(_14018_),
    .B2(_15046_),
    .ZN(_00908_));
 AOI21_X2 _23857_ (.A(_13998_),
    .B1(_14047_),
    .B2(_13952_),
    .ZN(_00909_));
 AOI21_X2 _23858_ (.A(_00908_),
    .B1(_00909_),
    .B2(_13951_),
    .ZN(_00910_));
 OAI21_X4 _23859_ (.A(_14156_),
    .B1(_14036_),
    .B2(_14014_),
    .ZN(_00911_));
 OAI21_X2 _23860_ (.A(_14112_),
    .B1(_00911_),
    .B2(_14021_),
    .ZN(_00912_));
 AOI21_X2 _23861_ (.A(_00910_),
    .B1(_00912_),
    .B2(_14012_),
    .ZN(_00913_));
 AOI221_X1 _23862_ (.A(_00773_),
    .B1(_00904_),
    .B2(_00907_),
    .C1(_00913_),
    .C2(_14034_),
    .ZN(_00914_));
 NOR3_X1 _23863_ (.A1(_14047_),
    .A2(_14078_),
    .A3(_00730_),
    .ZN(_00915_));
 OAI21_X1 _23864_ (.A(_13999_),
    .B1(_14176_),
    .B2(_14006_),
    .ZN(_00916_));
 OAI21_X1 _23865_ (.A(_14065_),
    .B1(_00915_),
    .B2(_00916_),
    .ZN(_00917_));
 NOR2_X1 _23866_ (.A1(_13990_),
    .A2(_00761_),
    .ZN(_00918_));
 AOI21_X1 _23867_ (.A(_13923_),
    .B1(_00850_),
    .B2(_00918_),
    .ZN(_00919_));
 NOR2_X1 _23868_ (.A1(_15020_),
    .A2(_13877_),
    .ZN(_00920_));
 AOI21_X1 _23869_ (.A(_14053_),
    .B1(_13966_),
    .B2(net1185),
    .ZN(_00921_));
 AOI21_X1 _23870_ (.A(_00920_),
    .B1(_00921_),
    .B2(_13965_),
    .ZN(_00922_));
 AND2_X1 _23871_ (.A1(_13877_),
    .A2(_00653_),
    .ZN(_00923_));
 AOI22_X1 _23872_ (.A1(_14156_),
    .A2(_00840_),
    .B1(_00923_),
    .B2(_14079_),
    .ZN(_00924_));
 MUX2_X1 _23873_ (.A(_00922_),
    .B(_00924_),
    .S(_13990_),
    .Z(_00925_));
 AOI221_X1 _23874_ (.A(_00749_),
    .B1(_00917_),
    .B2(_00919_),
    .C1(_00925_),
    .C2(_14051_),
    .ZN(_00926_));
 AOI221_X2 _23875_ (.A(_13990_),
    .B1(_14004_),
    .B2(_13985_),
    .C1(_14021_),
    .C2(_13923_),
    .ZN(_00927_));
 NOR3_X1 _23876_ (.A1(_14039_),
    .A2(_13924_),
    .A3(_14099_),
    .ZN(_00928_));
 OAI21_X1 _23877_ (.A(_13960_),
    .B1(_13964_),
    .B2(_14039_),
    .ZN(_00929_));
 AOI21_X1 _23878_ (.A(_00928_),
    .B1(_00929_),
    .B2(_15027_),
    .ZN(_00930_));
 OAI21_X1 _23879_ (.A(_00927_),
    .B1(_00930_),
    .B2(net1115),
    .ZN(_00931_));
 OAI21_X1 _23880_ (.A(_14029_),
    .B1(_13984_),
    .B2(_14151_),
    .ZN(_00932_));
 AOI21_X1 _23881_ (.A(_14031_),
    .B1(_14068_),
    .B2(_00932_),
    .ZN(_00933_));
 AOI21_X1 _23882_ (.A(_14003_),
    .B1(_14026_),
    .B2(_14039_),
    .ZN(_00934_));
 AOI21_X1 _23883_ (.A(_14089_),
    .B1(_14113_),
    .B2(_15018_),
    .ZN(_00935_));
 OAI22_X1 _23884_ (.A1(_14029_),
    .A2(_00934_),
    .B1(_00935_),
    .B2(_14051_),
    .ZN(_00936_));
 OAI21_X1 _23885_ (.A(_13992_),
    .B1(_00933_),
    .B2(_00936_),
    .ZN(_00937_));
 AOI21_X1 _23886_ (.A(_14105_),
    .B1(_00931_),
    .B2(_00937_),
    .ZN(_00938_));
 OR4_X2 _23887_ (.A1(_00926_),
    .A2(_00914_),
    .A3(_00902_),
    .A4(_00938_),
    .ZN(_00095_));
 XOR2_X2 _23888_ (.A(\sa00_sr[1] ),
    .B(_08987_),
    .Z(_00939_));
 XNOR2_X2 _23889_ (.A(_09153_),
    .B(_00939_),
    .ZN(_00940_));
 XOR2_X2 _23890_ (.A(net1104),
    .B(net919),
    .Z(_00941_));
 XNOR2_X2 _23891_ (.A(net631),
    .B(_00941_),
    .ZN(_00942_));
 XNOR2_X2 _23892_ (.A(_00940_),
    .B(_00942_),
    .ZN(_00943_));
 MUX2_X2 _23893_ (.A(_00464_),
    .B(_00943_),
    .S(_09195_),
    .Z(_00944_));
 XOR2_X2 _23894_ (.A(_06465_),
    .B(_00944_),
    .Z(_00945_));
 INV_X8 _23895_ (.A(net835),
    .ZN(_00946_));
 BUF_X4 clone288 (.A(net843),
    .Z(net836));
 BUF_X8 clone417 (.A(_00961_),
    .Z(net945));
 XNOR2_X1 _23898_ (.A(_08986_),
    .B(net691),
    .ZN(_00948_));
 NAND3_X4 _23899_ (.A1(_06450_),
    .A2(_09118_),
    .A3(net946),
    .ZN(_00949_));
 OR3_X1 _23900_ (.A1(_06450_),
    .A2(_11841_),
    .A3(_09153_),
    .ZN(_00950_));
 AOI21_X4 _23901_ (.A(_00948_),
    .B1(_00950_),
    .B2(_00949_),
    .ZN(_00951_));
 XOR2_X1 _23902_ (.A(_08986_),
    .B(net691),
    .Z(_00952_));
 INV_X1 _23903_ (.A(_06450_),
    .ZN(_00953_));
 NAND3_X1 _23904_ (.A1(_00953_),
    .A2(_09116_),
    .A3(_09153_),
    .ZN(_00954_));
 OR3_X1 _23905_ (.A1(_00953_),
    .A2(_09030_),
    .A3(_09153_),
    .ZN(_00955_));
 AOI21_X1 _23906_ (.A(_00952_),
    .B1(_00954_),
    .B2(_00955_),
    .ZN(_00956_));
 NAND3_X2 _23907_ (.A1(_00953_),
    .A2(_09179_),
    .A3(_00465_),
    .ZN(_00957_));
 NAND2_X1 _23908_ (.A1(_06450_),
    .A2(_09179_),
    .ZN(_00958_));
 OAI21_X2 _23909_ (.A(_00957_),
    .B1(_00958_),
    .B2(_00465_),
    .ZN(_00959_));
 OR3_X4 _23910_ (.A1(_00951_),
    .A2(_00956_),
    .A3(_00959_),
    .ZN(_00960_));
 INV_X8 _23911_ (.A(_00960_),
    .ZN(_00961_));
 BUF_X16 _23912_ (.A(_00961_),
    .Z(_00962_));
 BUF_X32 _23913_ (.A(_00962_),
    .Z(_15061_));
 XOR2_X2 _23914_ (.A(net694),
    .B(_09040_),
    .Z(_00963_));
 XOR2_X1 _23915_ (.A(_08987_),
    .B(_00963_),
    .Z(_00964_));
 NAND3_X1 _23916_ (.A1(_06480_),
    .A2(_09116_),
    .A3(_11882_),
    .ZN(_00965_));
 NOR2_X1 _23917_ (.A1(_06480_),
    .A2(_09028_),
    .ZN(_00966_));
 NAND2_X1 _23918_ (.A1(_11875_),
    .A2(_00966_),
    .ZN(_00967_));
 AOI21_X2 _23919_ (.A(_00964_),
    .B1(_00965_),
    .B2(_00967_),
    .ZN(_00968_));
 XNOR2_X1 _23920_ (.A(_08987_),
    .B(_00963_),
    .ZN(_00969_));
 NAND2_X1 _23921_ (.A1(_11882_),
    .A2(_00966_),
    .ZN(_00970_));
 NAND3_X1 _23922_ (.A1(_06480_),
    .A2(_09075_),
    .A3(_11875_),
    .ZN(_00971_));
 AOI21_X2 _23923_ (.A(_00969_),
    .B1(_00970_),
    .B2(_00971_),
    .ZN(_00972_));
 INV_X1 _23924_ (.A(_06480_),
    .ZN(_00973_));
 NAND3_X1 _23925_ (.A1(_00973_),
    .A2(_09730_),
    .A3(_00466_),
    .ZN(_00974_));
 NAND2_X1 _23926_ (.A1(_06480_),
    .A2(_09730_),
    .ZN(_00975_));
 OAI21_X2 _23927_ (.A(_00974_),
    .B1(_00975_),
    .B2(_00466_),
    .ZN(_00976_));
 NOR3_X4 _23928_ (.A1(_00976_),
    .A2(_00972_),
    .A3(_00968_),
    .ZN(_00977_));
 INV_X4 _23929_ (.A(net937),
    .ZN(_00978_));
 BUF_X8 _23930_ (.A(_00978_),
    .Z(_00979_));
 BUF_X4 _23931_ (.A(_00979_),
    .Z(_00980_));
 BUF_X8 _23932_ (.A(_00980_),
    .Z(_00981_));
 BUF_X8 _23933_ (.A(_00981_),
    .Z(_15077_));
 BUF_X1 rebuffer298 (.A(_00945_),
    .Z(net843));
 BUF_X4 _23935_ (.A(net940),
    .Z(_00982_));
 BUF_X4 _23936_ (.A(_00982_),
    .Z(_00983_));
 BUF_X4 _23937_ (.A(_00983_),
    .Z(_15070_));
 XNOR2_X1 _23938_ (.A(_09071_),
    .B(_09152_),
    .ZN(_00984_));
 XNOR2_X1 _23939_ (.A(_09014_),
    .B(_00984_),
    .ZN(_00985_));
 XNOR2_X1 _23940_ (.A(_09067_),
    .B(_00985_),
    .ZN(_00986_));
 MUX2_X1 _23941_ (.A(\text_in_r[111] ),
    .B(_00986_),
    .S(_09175_),
    .Z(_00987_));
 XNOR2_X2 _23942_ (.A(_06564_),
    .B(_00987_),
    .ZN(_00988_));
 INV_X2 _23943_ (.A(_00988_),
    .ZN(_00989_));
 INV_X1 _23944_ (.A(_06542_),
    .ZN(_00990_));
 BUF_X8 _23945_ (.A(_08994_),
    .Z(_00991_));
 XNOR2_X1 _23946_ (.A(_09187_),
    .B(_09166_),
    .ZN(_00992_));
 NOR3_X1 _23947_ (.A1(_00990_),
    .A2(_00991_),
    .A3(_00992_),
    .ZN(_00993_));
 NOR3_X1 _23948_ (.A1(_06542_),
    .A2(_00991_),
    .A3(_00992_),
    .ZN(_00994_));
 XNOR2_X1 _23949_ (.A(_09070_),
    .B(_09065_),
    .ZN(_00995_));
 XNOR2_X2 _23950_ (.A(_09190_),
    .B(_00995_),
    .ZN(_00996_));
 MUX2_X1 _23951_ (.A(_00993_),
    .B(_00994_),
    .S(_00996_),
    .Z(_00997_));
 XOR2_X1 _23952_ (.A(_09187_),
    .B(_09166_),
    .Z(_00998_));
 NOR3_X1 _23953_ (.A1(_06542_),
    .A2(_09103_),
    .A3(_00998_),
    .ZN(_00999_));
 NOR3_X1 _23954_ (.A1(_00990_),
    .A2(_09103_),
    .A3(_00998_),
    .ZN(_01000_));
 MUX2_X1 _23955_ (.A(_00999_),
    .B(_01000_),
    .S(_00996_),
    .Z(_01001_));
 NAND3_X1 _23956_ (.A1(_06542_),
    .A2(_09180_),
    .A3(\text_in_r[109] ),
    .ZN(_01002_));
 NAND2_X1 _23957_ (.A1(_00990_),
    .A2(_09180_),
    .ZN(_01003_));
 OAI21_X2 _23958_ (.A(_01002_),
    .B1(_01003_),
    .B2(\text_in_r[109] ),
    .ZN(_01004_));
 OR3_X2 _23959_ (.A1(_00997_),
    .A2(_01001_),
    .A3(_01004_),
    .ZN(_01005_));
 BUF_X4 _23960_ (.A(_01005_),
    .Z(_01006_));
 CLKBUF_X3 _23961_ (.A(_01006_),
    .Z(_01007_));
 XNOR2_X1 _23962_ (.A(_09169_),
    .B(_11897_),
    .ZN(_01008_));
 XNOR2_X1 _23963_ (.A(_09066_),
    .B(_01008_),
    .ZN(_01009_));
 MUX2_X2 _23964_ (.A(\text_in_r[110] ),
    .B(_01009_),
    .S(net951),
    .Z(_01010_));
 XOR2_X2 _23965_ (.A(_06555_),
    .B(_01010_),
    .Z(_01011_));
 NAND2_X1 _23966_ (.A1(_06527_),
    .A2(_09175_),
    .ZN(_01012_));
 INV_X1 _23967_ (.A(_06527_),
    .ZN(_01013_));
 NAND2_X1 _23968_ (.A1(_01013_),
    .A2(_09175_),
    .ZN(_01014_));
 XNOR2_X1 _23969_ (.A(_09094_),
    .B(_09152_),
    .ZN(_01015_));
 XNOR2_X2 _23970_ (.A(_09163_),
    .B(_01015_),
    .ZN(_01016_));
 XNOR2_X1 _23971_ (.A(_11907_),
    .B(_01016_),
    .ZN(_01017_));
 MUX2_X2 _23972_ (.A(_01012_),
    .B(_01014_),
    .S(_01017_),
    .Z(_01018_));
 NOR3_X2 _23973_ (.A1(_01013_),
    .A2(_09138_),
    .A3(\text_in_r[108] ),
    .ZN(_01019_));
 NOR2_X1 _23974_ (.A1(_06527_),
    .A2(_10571_),
    .ZN(_01020_));
 AOI21_X4 _23975_ (.A(_01019_),
    .B1(_01020_),
    .B2(\text_in_r[108] ),
    .ZN(_01021_));
 NAND2_X1 _23976_ (.A1(_01018_),
    .A2(_01021_),
    .ZN(_01022_));
 BUF_X4 _23977_ (.A(_01022_),
    .Z(_01023_));
 BUF_X4 _23978_ (.A(_01023_),
    .Z(_01024_));
 NOR2_X2 _23979_ (.A1(_01011_),
    .A2(_01024_),
    .ZN(_01025_));
 BUF_X4 _23980_ (.A(_00979_),
    .Z(_01026_));
 BUF_X4 _23981_ (.A(_01026_),
    .Z(_01027_));
 BUF_X1 split188 (.A(_15270_),
    .Z(net188));
 INV_X1 _23983_ (.A(_06510_),
    .ZN(_01029_));
 NOR2_X1 _23984_ (.A1(_01029_),
    .A2(_08995_),
    .ZN(_01030_));
 NOR2_X1 _23985_ (.A1(_06510_),
    .A2(_08995_),
    .ZN(_01031_));
 XNOR2_X1 _23986_ (.A(_09186_),
    .B(_09152_),
    .ZN(_01032_));
 XNOR2_X2 _23987_ (.A(_09037_),
    .B(_09092_),
    .ZN(_01033_));
 XNOR2_X2 _23988_ (.A(_01032_),
    .B(_01033_),
    .ZN(_01034_));
 XNOR2_X1 _23989_ (.A(_09094_),
    .B(_09151_),
    .ZN(_01035_));
 XNOR2_X1 _23990_ (.A(_09041_),
    .B(_01035_),
    .ZN(_01036_));
 XNOR2_X2 _23991_ (.A(_01034_),
    .B(_01036_),
    .ZN(_01037_));
 MUX2_X2 _23992_ (.A(_01030_),
    .B(_01031_),
    .S(_01037_),
    .Z(_01038_));
 BUF_X8 _23993_ (.A(_01038_),
    .Z(_01039_));
 BUF_X4 _23994_ (.A(_01039_),
    .Z(_01040_));
 OR3_X2 _23995_ (.A1(_01029_),
    .A2(_09075_),
    .A3(\text_in_r[107] ),
    .ZN(_01041_));
 NAND3_X2 _23996_ (.A1(_01029_),
    .A2(_08995_),
    .A3(\text_in_r[107] ),
    .ZN(_01042_));
 NAND2_X4 _23997_ (.A1(_01041_),
    .A2(_01042_),
    .ZN(_01043_));
 BUF_X8 _23998_ (.A(_01043_),
    .Z(_01044_));
 BUF_X4 _23999_ (.A(_01044_),
    .Z(_01045_));
 NOR3_X2 _24000_ (.A1(net1032),
    .A2(_01040_),
    .A3(_01045_),
    .ZN(_01046_));
 BUF_X4 _24001_ (.A(_15052_),
    .Z(_01047_));
 NAND2_X1 _24002_ (.A1(_06510_),
    .A2(net951),
    .ZN(_01048_));
 NAND2_X1 _24003_ (.A1(_01029_),
    .A2(net951),
    .ZN(_01049_));
 MUX2_X2 _24004_ (.A(_01048_),
    .B(_01049_),
    .S(_01037_),
    .Z(_01050_));
 BUF_X8 _24005_ (.A(_01050_),
    .Z(_01051_));
 BUF_X4 _24006_ (.A(_01051_),
    .Z(_01052_));
 AND2_X1 _24007_ (.A1(_01041_),
    .A2(_01042_),
    .ZN(_01053_));
 BUF_X8 _24008_ (.A(_01053_),
    .Z(_01054_));
 BUF_X8 _24009_ (.A(_01054_),
    .Z(_01055_));
 AOI21_X1 _24010_ (.A(_01047_),
    .B1(_01052_),
    .B2(_01055_),
    .ZN(_01056_));
 NOR3_X1 _24011_ (.A1(_01027_),
    .A2(_01046_),
    .A3(_01056_),
    .ZN(_01057_));
 AOI21_X4 _24012_ (.A(_00960_),
    .B1(_01052_),
    .B2(_01055_),
    .ZN(_01058_));
 BUF_X8 _24013_ (.A(_15054_),
    .Z(_01059_));
 NOR2_X4 _24014_ (.A1(_15059_),
    .A2(_01059_),
    .ZN(_01060_));
 NOR3_X2 _24015_ (.A1(_01040_),
    .A2(_01045_),
    .A3(_01060_),
    .ZN(_01061_));
 NOR3_X1 _24016_ (.A1(_00983_),
    .A2(_01058_),
    .A3(_01061_),
    .ZN(_01062_));
 OAI21_X1 _24017_ (.A(_01025_),
    .B1(_01057_),
    .B2(_01062_),
    .ZN(_01063_));
 CLKBUF_X3 _24018_ (.A(_01011_),
    .Z(_01064_));
 AND2_X1 _24019_ (.A1(_01018_),
    .A2(_01021_),
    .ZN(_01065_));
 BUF_X4 _24020_ (.A(_01065_),
    .Z(_01066_));
 BUF_X4 _24021_ (.A(_01066_),
    .Z(_01067_));
 BUF_X4 _24022_ (.A(_01067_),
    .Z(_01068_));
 BUF_X1 rebuffer407 (.A(_09319_),
    .Z(net870));
 INV_X2 _24024_ (.A(net1033),
    .ZN(_01070_));
 AOI21_X4 _24025_ (.A(_00978_),
    .B1(_01051_),
    .B2(_01054_),
    .ZN(_01071_));
 NAND2_X1 _24026_ (.A1(_01070_),
    .A2(_01071_),
    .ZN(_01072_));
 BUF_X8 _24027_ (.A(_15059_),
    .Z(_01073_));
 INV_X4 _24028_ (.A(_01073_),
    .ZN(_01074_));
 NOR3_X4 _24029_ (.A1(_01074_),
    .A2(_01040_),
    .A3(_01045_),
    .ZN(_01075_));
 OAI21_X1 _24030_ (.A(_01027_),
    .B1(_01058_),
    .B2(_01075_),
    .ZN(_01076_));
 NAND4_X1 _24031_ (.A1(_01064_),
    .A2(_01068_),
    .A3(_01072_),
    .A4(_01076_),
    .ZN(_01077_));
 AND4_X1 _24032_ (.A1(_00989_),
    .A2(_01007_),
    .A3(_01063_),
    .A4(_01077_),
    .ZN(_01078_));
 NAND2_X2 _24033_ (.A1(_01050_),
    .A2(_01053_),
    .ZN(_01079_));
 BUF_X4 _24034_ (.A(_01079_),
    .Z(_01080_));
 BUF_X4 _24035_ (.A(_01080_),
    .Z(_01081_));
 NOR3_X2 _24036_ (.A1(net937),
    .A2(_01039_),
    .A3(_01044_),
    .ZN(_01082_));
 BUF_X4 _24037_ (.A(_01082_),
    .Z(_01083_));
 BUF_X8 _24038_ (.A(net687),
    .Z(_01084_));
 AOI221_X2 _24039_ (.A(_01011_),
    .B1(_01081_),
    .B2(_15075_),
    .C1(_01083_),
    .C2(net682),
    .ZN(_01085_));
 AOI21_X4 _24040_ (.A(_01084_),
    .B1(_01051_),
    .B2(_01054_),
    .ZN(_01086_));
 BUF_X8 _24041_ (.A(_15064_),
    .Z(_01087_));
 NOR3_X2 _24042_ (.A1(_01087_),
    .A2(_01040_),
    .A3(_01045_),
    .ZN(_01088_));
 OAI21_X1 _24043_ (.A(_15070_),
    .B1(_01086_),
    .B2(_01088_),
    .ZN(_01089_));
 NOR2_X4 _24044_ (.A1(_01038_),
    .A2(_01043_),
    .ZN(_01090_));
 BUF_X4 _24045_ (.A(_01090_),
    .Z(_01091_));
 NAND2_X4 _24046_ (.A1(_00979_),
    .A2(_01091_),
    .ZN(_01092_));
 OAI21_X1 _24047_ (.A(_01089_),
    .B1(_01092_),
    .B2(_01073_),
    .ZN(_01093_));
 AOI21_X1 _24048_ (.A(_01085_),
    .B1(_01093_),
    .B2(_01064_),
    .ZN(_01094_));
 NAND2_X1 _24049_ (.A1(_00988_),
    .A2(_01007_),
    .ZN(_01095_));
 BUF_X4 _24050_ (.A(_01024_),
    .Z(_01096_));
 NOR2_X2 _24051_ (.A1(_01059_),
    .A2(_00978_),
    .ZN(_01097_));
 AOI211_X2 _24052_ (.A(_01079_),
    .B(_01097_),
    .C1(net740),
    .C2(_00979_),
    .ZN(_01098_));
 BUF_X4 _24053_ (.A(_01090_),
    .Z(_01099_));
 BUF_X8 _24054_ (.A(net941),
    .Z(_15050_));
 MUX2_X1 _24055_ (.A(_15066_),
    .B(_15050_),
    .S(_00978_),
    .Z(_01100_));
 OAI21_X1 _24056_ (.A(_01011_),
    .B1(_01099_),
    .B2(_01100_),
    .ZN(_01101_));
 NOR3_X1 _24057_ (.A1(_01096_),
    .A2(_01098_),
    .A3(_01101_),
    .ZN(_01102_));
 BUF_X4 _24058_ (.A(_15062_),
    .Z(_01103_));
 NAND2_X1 _24059_ (.A1(_01103_),
    .A2(_01083_),
    .ZN(_01104_));
 AOI21_X4 _24060_ (.A(net940),
    .B1(_01052_),
    .B2(_01055_),
    .ZN(_01105_));
 NOR3_X4 _24061_ (.A1(_00978_),
    .A2(_01039_),
    .A3(_01044_),
    .ZN(_01106_));
 NOR2_X2 _24062_ (.A1(_01105_),
    .A2(_01106_),
    .ZN(_01107_));
 INV_X2 _24063_ (.A(_01047_),
    .ZN(_01108_));
 OAI21_X4 _24064_ (.A(_00982_),
    .B1(_01040_),
    .B2(_01045_),
    .ZN(_01109_));
 OAI221_X2 _24065_ (.A(_01104_),
    .B1(_01107_),
    .B2(_01108_),
    .C1(_01109_),
    .C2(net682),
    .ZN(_01110_));
 AOI211_X2 _24066_ (.A(_01095_),
    .B(_01102_),
    .C1(_01110_),
    .C2(_01025_),
    .ZN(_01111_));
 NOR3_X1 _24067_ (.A1(_00983_),
    .A2(_01058_),
    .A3(_01046_),
    .ZN(_01112_));
 BUF_X8 _24068_ (.A(_15068_),
    .Z(_01113_));
 OAI21_X1 _24069_ (.A(_01113_),
    .B1(_01039_),
    .B2(_01044_),
    .ZN(_01114_));
 AND2_X1 _24070_ (.A1(_00983_),
    .A2(_01114_),
    .ZN(_01115_));
 NAND2_X1 _24071_ (.A1(net742),
    .A2(_01099_),
    .ZN(_01116_));
 AOI21_X1 _24072_ (.A(_01112_),
    .B1(_01115_),
    .B2(_01116_),
    .ZN(_01117_));
 INV_X8 _24073_ (.A(net687),
    .ZN(_01118_));
 NOR3_X4 _24074_ (.A1(_01118_),
    .A2(_01039_),
    .A3(_01044_),
    .ZN(_01119_));
 OAI21_X1 _24075_ (.A(_01119_),
    .B1(_00983_),
    .B2(net742),
    .ZN(_01120_));
 NAND2_X1 _24076_ (.A1(_01118_),
    .A2(_00981_),
    .ZN(_01121_));
 BUF_X4 _24077_ (.A(_01080_),
    .Z(_01122_));
 NOR2_X2 _24078_ (.A1(net844),
    .A2(_01122_),
    .ZN(_01123_));
 OAI21_X1 _24079_ (.A(_01120_),
    .B1(_01121_),
    .B2(_01123_),
    .ZN(_01124_));
 XNOR2_X2 _24080_ (.A(_06555_),
    .B(_01010_),
    .ZN(_01125_));
 MUX2_X1 _24081_ (.A(_01117_),
    .B(_01124_),
    .S(_01125_),
    .Z(_01126_));
 AOI22_X1 _24082_ (.A1(_01078_),
    .A2(_01094_),
    .B1(_01111_),
    .B2(_01126_),
    .ZN(_01127_));
 NOR2_X1 _24083_ (.A1(_01078_),
    .A2(_01111_),
    .ZN(_01128_));
 BUF_X4 _24084_ (.A(_01096_),
    .Z(_01129_));
 NAND2_X1 _24085_ (.A1(_01011_),
    .A2(_01022_),
    .ZN(_01130_));
 NAND3_X2 _24086_ (.A1(_01059_),
    .A2(_01051_),
    .A3(_01054_),
    .ZN(_01131_));
 AOI21_X1 _24087_ (.A(_00978_),
    .B1(_01079_),
    .B2(_01073_),
    .ZN(_01132_));
 AOI221_X1 _24088_ (.A(_01130_),
    .B1(_01131_),
    .B2(_01132_),
    .C1(_01083_),
    .C2(_01047_),
    .ZN(_01133_));
 OR2_X1 _24089_ (.A1(_00988_),
    .A2(_01133_),
    .ZN(_01134_));
 AOI21_X1 _24090_ (.A(_01046_),
    .B1(_01081_),
    .B2(net925),
    .ZN(_01135_));
 OAI22_X2 _24091_ (.A1(_01103_),
    .A2(_01092_),
    .B1(_01135_),
    .B2(_00981_),
    .ZN(_01136_));
 NOR2_X1 _24092_ (.A1(_01064_),
    .A2(_01068_),
    .ZN(_01137_));
 OR2_X1 _24093_ (.A1(_01026_),
    .A2(_01058_),
    .ZN(_01138_));
 AOI21_X4 _24094_ (.A(_01103_),
    .B1(_01052_),
    .B2(_01055_),
    .ZN(_01139_));
 NOR3_X4 _24095_ (.A1(_01043_),
    .A2(_01038_),
    .A3(net503),
    .ZN(_01140_));
 OR2_X2 _24096_ (.A1(_01139_),
    .A2(_01140_),
    .ZN(_01141_));
 BUF_X4 _24097_ (.A(net937),
    .Z(_01142_));
 BUF_X4 _24098_ (.A(_01142_),
    .Z(_01143_));
 CLKBUF_X3 _24099_ (.A(_01143_),
    .Z(_01144_));
 OAI221_X2 _24100_ (.A(_01064_),
    .B1(_01123_),
    .B2(_01138_),
    .C1(_01141_),
    .C2(_01144_),
    .ZN(_01145_));
 BUF_X4 _24101_ (.A(_01091_),
    .Z(_01146_));
 BUF_X4 _24102_ (.A(net923),
    .Z(_01147_));
 OAI21_X1 _24103_ (.A(_01131_),
    .B1(_01146_),
    .B2(_01147_),
    .ZN(_01148_));
 AOI22_X1 _24104_ (.A1(_01144_),
    .A2(_01148_),
    .B1(_01105_),
    .B2(net1056),
    .ZN(_01149_));
 OAI21_X2 _24105_ (.A(_01145_),
    .B1(_01149_),
    .B2(_01064_),
    .ZN(_01150_));
 BUF_X4 _24106_ (.A(_01068_),
    .Z(_01151_));
 AOI221_X2 _24107_ (.A(_01134_),
    .B1(_01136_),
    .B2(_01137_),
    .C1(_01150_),
    .C2(_01151_),
    .ZN(_01152_));
 NOR3_X4 _24108_ (.A1(_00997_),
    .A2(_01001_),
    .A3(_01004_),
    .ZN(_01153_));
 BUF_X4 _24109_ (.A(_01153_),
    .Z(_01154_));
 BUF_X4 _24110_ (.A(_01154_),
    .Z(_01155_));
 BUF_X4 _24111_ (.A(_01155_),
    .Z(_01156_));
 NAND2_X1 _24112_ (.A1(_00988_),
    .A2(_01129_),
    .ZN(_01157_));
 BUF_X4 _24113_ (.A(_01080_),
    .Z(_01158_));
 CLKBUF_X3 _24114_ (.A(_01158_),
    .Z(_01159_));
 NAND2_X2 _24115_ (.A1(_00961_),
    .A2(_01142_),
    .ZN(_01160_));
 OAI21_X1 _24116_ (.A(_01160_),
    .B1(_00962_),
    .B2(net1030),
    .ZN(_01161_));
 XNOR2_X1 _24117_ (.A(_01159_),
    .B(_01161_),
    .ZN(_01162_));
 OAI21_X4 _24118_ (.A(_01084_),
    .B1(_01040_),
    .B2(_01045_),
    .ZN(_01163_));
 NAND3_X4 _24119_ (.A1(_00961_),
    .A2(_01051_),
    .A3(_01054_),
    .ZN(_01164_));
 AND3_X4 _24120_ (.A1(_01163_),
    .A2(_00982_),
    .A3(_01164_),
    .ZN(_01165_));
 NAND3_X4 _24121_ (.A1(_01054_),
    .A2(_01051_),
    .A3(net1032),
    .ZN(_01166_));
 OAI21_X1 _24122_ (.A(_01166_),
    .B1(_01091_),
    .B2(_01113_),
    .ZN(_01167_));
 AOI21_X1 _24123_ (.A(_01165_),
    .B1(_01167_),
    .B2(_00981_),
    .ZN(_01168_));
 MUX2_X1 _24124_ (.A(_01162_),
    .B(_01168_),
    .S(_01064_),
    .Z(_01169_));
 BUF_X4 _24125_ (.A(_01096_),
    .Z(_01170_));
 BUF_X4 _24126_ (.A(_00978_),
    .Z(_01171_));
 BUF_X4 _24127_ (.A(_01171_),
    .Z(_01172_));
 NOR3_X1 _24128_ (.A1(_01172_),
    .A2(_01139_),
    .A3(_01119_),
    .ZN(_01173_));
 BUF_X4 _24129_ (.A(_00982_),
    .Z(_01174_));
 NOR3_X4 _24130_ (.A1(net1033),
    .A2(_01040_),
    .A3(_01045_),
    .ZN(_01175_));
 NOR3_X1 _24131_ (.A1(_01175_),
    .A2(_01056_),
    .A3(_01174_),
    .ZN(_01176_));
 NOR3_X1 _24132_ (.A1(_01064_),
    .A2(_01173_),
    .A3(_01176_),
    .ZN(_01177_));
 OAI21_X2 _24133_ (.A(_15057_),
    .B1(_01039_),
    .B2(_01044_),
    .ZN(_01178_));
 OAI21_X1 _24134_ (.A(_01178_),
    .B1(_01080_),
    .B2(_00961_),
    .ZN(_01179_));
 AOI221_X2 _24135_ (.A(_01125_),
    .B1(_01179_),
    .B2(_01171_),
    .C1(_01071_),
    .C2(_01074_),
    .ZN(_01180_));
 OR3_X1 _24136_ (.A1(_01170_),
    .A2(_01177_),
    .A3(_01180_),
    .ZN(_01181_));
 OAI221_X2 _24137_ (.A(_01156_),
    .B1(_01169_),
    .B2(_01157_),
    .C1(_00989_),
    .C2(_01181_),
    .ZN(_01182_));
 OAI221_X1 _24138_ (.A(_01127_),
    .B1(_01128_),
    .B2(_01129_),
    .C1(_01182_),
    .C2(_01152_),
    .ZN(_00096_));
 NOR2_X2 _24139_ (.A1(_00989_),
    .A2(_01125_),
    .ZN(_01183_));
 NAND2_X4 _24140_ (.A1(_01023_),
    .A2(_01154_),
    .ZN(_01184_));
 CLKBUF_X3 _24141_ (.A(_01172_),
    .Z(_01185_));
 OAI21_X1 _24142_ (.A(_01108_),
    .B1(_01040_),
    .B2(_01045_),
    .ZN(_01186_));
 AOI21_X1 _24143_ (.A(_01185_),
    .B1(_01131_),
    .B2(_01186_),
    .ZN(_01187_));
 AOI21_X1 _24144_ (.A(_01142_),
    .B1(_01163_),
    .B2(_01164_),
    .ZN(_01188_));
 OR2_X1 _24145_ (.A1(_01187_),
    .A2(_01188_),
    .ZN(_01189_));
 CLKBUF_X3 _24146_ (.A(_01007_),
    .Z(_01190_));
 CLKBUF_X3 _24147_ (.A(_01146_),
    .Z(_01191_));
 BUF_X4 _24148_ (.A(_15066_),
    .Z(_01192_));
 AOI21_X1 _24149_ (.A(net743),
    .B1(_01191_),
    .B2(_01192_),
    .ZN(_01193_));
 OAI221_X1 _24150_ (.A(_01190_),
    .B1(_01193_),
    .B2(_15077_),
    .C1(_01092_),
    .C2(net950),
    .ZN(_01194_));
 NOR2_X1 _24151_ (.A1(_01129_),
    .A2(_01194_),
    .ZN(_01195_));
 NOR3_X4 _24152_ (.A1(_00960_),
    .A2(_01038_),
    .A3(_01043_),
    .ZN(_01196_));
 AOI21_X4 _24153_ (.A(_01073_),
    .B1(_01051_),
    .B2(_01054_),
    .ZN(_01197_));
 NOR3_X1 _24154_ (.A1(_01172_),
    .A2(_01196_),
    .A3(_01197_),
    .ZN(_01198_));
 MUX2_X1 _24155_ (.A(_01108_),
    .B(net741),
    .S(_01159_),
    .Z(_01199_));
 AOI21_X1 _24156_ (.A(_01198_),
    .B1(_01199_),
    .B2(_15077_),
    .ZN(_01200_));
 OAI21_X2 _24157_ (.A(_01118_),
    .B1(_01039_),
    .B2(_01044_),
    .ZN(_01201_));
 NAND3_X1 _24158_ (.A1(_01113_),
    .A2(_01052_),
    .A3(_01055_),
    .ZN(_01202_));
 AOI21_X1 _24159_ (.A(_01185_),
    .B1(_01201_),
    .B2(_01202_),
    .ZN(_01203_));
 OAI21_X1 _24160_ (.A(_01070_),
    .B1(_01040_),
    .B2(_01045_),
    .ZN(_01204_));
 AOI21_X1 _24161_ (.A(_01144_),
    .B1(_01131_),
    .B2(_01204_),
    .ZN(_01205_));
 OAI21_X1 _24162_ (.A(_01170_),
    .B1(_01203_),
    .B2(_01205_),
    .ZN(_01206_));
 AOI22_X1 _24163_ (.A1(_01151_),
    .A2(_01200_),
    .B1(_01206_),
    .B2(_01190_),
    .ZN(_01207_));
 OAI221_X1 _24164_ (.A(_01183_),
    .B1(_01184_),
    .B2(_01189_),
    .C1(_01195_),
    .C2(_01207_),
    .ZN(_01208_));
 NOR2_X2 _24165_ (.A1(_00988_),
    .A2(_01125_),
    .ZN(_01209_));
 OAI21_X4 _24166_ (.A(_00979_),
    .B1(_01040_),
    .B2(_01045_),
    .ZN(_01210_));
 INV_X4 _24167_ (.A(_01113_),
    .ZN(_01211_));
 BUF_X4 _24168_ (.A(net835),
    .Z(_01212_));
 NOR2_X2 _24169_ (.A1(_01212_),
    .A2(_01099_),
    .ZN(_01213_));
 NOR2_X1 _24170_ (.A1(_01175_),
    .A2(_01213_),
    .ZN(_01214_));
 OAI221_X1 _24171_ (.A(_01129_),
    .B1(_01210_),
    .B2(_01211_),
    .C1(_01214_),
    .C2(_15077_),
    .ZN(_01215_));
 NOR2_X1 _24172_ (.A1(net737),
    .A2(_01075_),
    .ZN(_01216_));
 OAI221_X1 _24173_ (.A(_01151_),
    .B1(_01210_),
    .B2(_01192_),
    .C1(_01216_),
    .C2(_15077_),
    .ZN(_01217_));
 NAND4_X1 _24174_ (.A1(_01156_),
    .A2(_01209_),
    .A3(_01215_),
    .A4(_01217_),
    .ZN(_01218_));
 NOR2_X2 _24175_ (.A1(_00988_),
    .A2(_01011_),
    .ZN(_01219_));
 NAND2_X1 _24176_ (.A1(_01154_),
    .A2(_01219_),
    .ZN(_01220_));
 AOI21_X1 _24177_ (.A(_01023_),
    .B1(_01196_),
    .B2(net8),
    .ZN(_01221_));
 NOR2_X1 _24178_ (.A1(net1032),
    .A2(_01090_),
    .ZN(_01222_));
 NOR2_X2 _24179_ (.A1(net8),
    .A2(_01079_),
    .ZN(_01223_));
 OAI21_X1 _24180_ (.A(_01171_),
    .B1(_01222_),
    .B2(_01223_),
    .ZN(_01224_));
 AOI21_X4 _24181_ (.A(_00961_),
    .B1(_01051_),
    .B2(_01054_),
    .ZN(_01225_));
 OAI21_X1 _24182_ (.A(_01171_),
    .B1(_01196_),
    .B2(_01225_),
    .ZN(_01226_));
 NOR3_X4 _24183_ (.A1(net681),
    .A2(_01038_),
    .A3(_01043_),
    .ZN(_01227_));
 NOR2_X4 _24184_ (.A1(net738),
    .A2(net743),
    .ZN(_01228_));
 OAI21_X4 _24185_ (.A(_01226_),
    .B1(_01171_),
    .B2(_01228_),
    .ZN(_01229_));
 AOI221_X2 _24186_ (.A(_01220_),
    .B1(_01221_),
    .B2(_01224_),
    .C1(_01229_),
    .C2(_01024_),
    .ZN(_01230_));
 NAND2_X2 _24187_ (.A1(net1030),
    .A2(net938),
    .ZN(_01231_));
 AOI21_X1 _24188_ (.A(_01079_),
    .B1(_00978_),
    .B2(_01074_),
    .ZN(_01232_));
 INV_X1 _24189_ (.A(_15082_),
    .ZN(_01233_));
 AOI221_X2 _24190_ (.A(_01066_),
    .B1(_01232_),
    .B2(_01231_),
    .C1(_01122_),
    .C2(_01233_),
    .ZN(_01234_));
 OR2_X1 _24191_ (.A1(_01086_),
    .A2(_01227_),
    .ZN(_01235_));
 MUX2_X1 _24192_ (.A(_01167_),
    .B(_01235_),
    .S(_00980_),
    .Z(_01236_));
 AOI21_X2 _24193_ (.A(_01234_),
    .B1(_01236_),
    .B2(_01068_),
    .ZN(_01237_));
 NAND2_X1 _24194_ (.A1(_00989_),
    .A2(_01125_),
    .ZN(_01238_));
 NOR2_X1 _24195_ (.A1(_01155_),
    .A2(_01238_),
    .ZN(_01239_));
 NOR2_X2 _24196_ (.A1(_00989_),
    .A2(_01011_),
    .ZN(_01240_));
 MUX2_X1 _24197_ (.A(_01103_),
    .B(_15066_),
    .S(net938),
    .Z(_01241_));
 BUF_X4 _24198_ (.A(_01006_),
    .Z(_01242_));
 NAND2_X1 _24199_ (.A1(_01081_),
    .A2(_01242_),
    .ZN(_01243_));
 OAI221_X1 _24200_ (.A(_01067_),
    .B1(_01081_),
    .B2(net686),
    .C1(_01243_),
    .C2(_15078_),
    .ZN(_01244_));
 NOR2_X1 _24201_ (.A1(_01067_),
    .A2(_01242_),
    .ZN(_01245_));
 NAND3_X4 _24202_ (.A1(_01047_),
    .A2(_01051_),
    .A3(_01054_),
    .ZN(_01246_));
 NAND3_X1 _24203_ (.A1(_01172_),
    .A2(_01178_),
    .A3(_01246_),
    .ZN(_01247_));
 AOI21_X4 _24204_ (.A(net1033),
    .B1(_01051_),
    .B2(_01054_),
    .ZN(_01248_));
 OAI21_X1 _24205_ (.A(_01174_),
    .B1(_01196_),
    .B2(_01248_),
    .ZN(_01249_));
 NAND3_X1 _24206_ (.A1(_01245_),
    .A2(_01247_),
    .A3(_01249_),
    .ZN(_01250_));
 AND3_X1 _24207_ (.A1(_01240_),
    .A2(_01244_),
    .A3(_01250_),
    .ZN(_01251_));
 NOR2_X2 _24208_ (.A1(_01067_),
    .A2(_01154_),
    .ZN(_01252_));
 XNOR2_X2 _24209_ (.A(net520),
    .B(_01090_),
    .ZN(_01253_));
 AOI21_X1 _24210_ (.A(_01198_),
    .B1(_01253_),
    .B2(_01185_),
    .ZN(_01254_));
 NAND2_X1 _24211_ (.A1(_01252_),
    .A2(_01254_),
    .ZN(_01255_));
 AOI221_X2 _24212_ (.A(_01230_),
    .B1(_01237_),
    .B2(_01239_),
    .C1(_01251_),
    .C2(_01255_),
    .ZN(_01256_));
 NAND3_X1 _24213_ (.A1(_00983_),
    .A2(_01163_),
    .A3(_01246_),
    .ZN(_01257_));
 BUF_X4 _24214_ (.A(_01081_),
    .Z(_01258_));
 AOI21_X1 _24215_ (.A(_01196_),
    .B1(_01258_),
    .B2(_01073_),
    .ZN(_01259_));
 OAI21_X1 _24216_ (.A(_01257_),
    .B1(_01259_),
    .B2(_15070_),
    .ZN(_01260_));
 NAND3_X2 _24217_ (.A1(_01142_),
    .A2(_01052_),
    .A3(_01055_),
    .ZN(_01261_));
 AOI21_X1 _24218_ (.A(net945),
    .B1(_01210_),
    .B2(_01261_),
    .ZN(_01262_));
 AOI221_X2 _24219_ (.A(_01262_),
    .B1(_01058_),
    .B2(_01212_),
    .C1(net682),
    .C2(_01083_),
    .ZN(_01263_));
 MUX2_X1 _24220_ (.A(_01260_),
    .B(_01263_),
    .S(_01151_),
    .Z(_01264_));
 NAND3_X1 _24221_ (.A1(_01190_),
    .A2(_01264_),
    .A3(_01209_),
    .ZN(_01265_));
 NAND4_X1 _24222_ (.A1(_01208_),
    .A2(_01256_),
    .A3(_01218_),
    .A4(_01265_),
    .ZN(_00097_));
 AND3_X1 _24223_ (.A1(_01018_),
    .A2(_01021_),
    .A3(_01006_),
    .ZN(_01266_));
 NAND3_X2 _24224_ (.A1(net942),
    .A2(_01052_),
    .A3(_01055_),
    .ZN(_01267_));
 NAND2_X1 _24225_ (.A1(_01143_),
    .A2(_01267_),
    .ZN(_01268_));
 OAI221_X2 _24226_ (.A(_01266_),
    .B1(_01268_),
    .B2(_01213_),
    .C1(_00983_),
    .C2(_01073_),
    .ZN(_01269_));
 OAI21_X4 _24227_ (.A(_15064_),
    .B1(_01039_),
    .B2(_01044_),
    .ZN(_01270_));
 AOI21_X1 _24228_ (.A(_00980_),
    .B1(_01270_),
    .B2(_01164_),
    .ZN(_01271_));
 NOR3_X4 _24229_ (.A1(_01113_),
    .A2(_01039_),
    .A3(_01044_),
    .ZN(_01272_));
 NOR2_X2 _24230_ (.A1(_00982_),
    .A2(_01272_),
    .ZN(_01273_));
 NAND2_X4 _24231_ (.A1(net740),
    .A2(_01080_),
    .ZN(_01274_));
 AOI21_X1 _24232_ (.A(_01271_),
    .B1(_01273_),
    .B2(_01274_),
    .ZN(_01275_));
 OAI211_X2 _24233_ (.A(_01183_),
    .B(_01269_),
    .C1(_01275_),
    .C2(_01184_),
    .ZN(_01276_));
 NOR3_X1 _24234_ (.A1(_01027_),
    .A2(_01088_),
    .A3(_01225_),
    .ZN(_01277_));
 NOR3_X1 _24235_ (.A1(_01174_),
    .A2(_01197_),
    .A3(_01272_),
    .ZN(_01278_));
 OAI21_X1 _24236_ (.A(_01252_),
    .B1(_01277_),
    .B2(_01278_),
    .ZN(_01279_));
 AND3_X2 _24237_ (.A1(_01171_),
    .A2(_01201_),
    .A3(_01267_),
    .ZN(_01280_));
 NAND2_X2 _24238_ (.A1(_01066_),
    .A2(_01153_),
    .ZN(_01281_));
 OR3_X4 _24239_ (.A1(_01165_),
    .A2(_01280_),
    .A3(_01281_),
    .ZN(_01282_));
 NAND2_X4 _24240_ (.A1(_01282_),
    .A2(_01279_),
    .ZN(_01283_));
 INV_X1 _24241_ (.A(_15057_),
    .ZN(_01284_));
 MUX2_X1 _24242_ (.A(_01073_),
    .B(_01284_),
    .S(_01142_),
    .Z(_01285_));
 OAI21_X4 _24243_ (.A(_01068_),
    .B1(_01146_),
    .B2(_01285_),
    .ZN(_01286_));
 NOR2_X2 _24244_ (.A1(_01118_),
    .A2(_01142_),
    .ZN(_01287_));
 OAI21_X1 _24245_ (.A(_01146_),
    .B1(_00980_),
    .B2(_01212_),
    .ZN(_01288_));
 OAI21_X1 _24246_ (.A(_01007_),
    .B1(_01287_),
    .B2(_01288_),
    .ZN(_01289_));
 AOI21_X2 _24247_ (.A(_01272_),
    .B1(_01158_),
    .B2(_01147_),
    .ZN(_01290_));
 NOR2_X4 _24248_ (.A1(net738),
    .A2(_00980_),
    .ZN(_01291_));
 AOI22_X4 _24249_ (.A1(_01027_),
    .A2(_01290_),
    .B1(_01291_),
    .B2(_01274_),
    .ZN(_01292_));
 NAND2_X2 _24250_ (.A1(_01023_),
    .A2(_01006_),
    .ZN(_01293_));
 OAI22_X4 _24251_ (.A1(_01286_),
    .A2(_01289_),
    .B1(_01293_),
    .B2(_01292_),
    .ZN(_01294_));
 NAND2_X1 _24252_ (.A1(_01192_),
    .A2(_01158_),
    .ZN(_01295_));
 AOI21_X1 _24253_ (.A(_01174_),
    .B1(_01166_),
    .B2(_01295_),
    .ZN(_01296_));
 NOR2_X1 _24254_ (.A1(_01023_),
    .A2(_01006_),
    .ZN(_01297_));
 OAI21_X1 _24255_ (.A(_01297_),
    .B1(_01109_),
    .B2(_01113_),
    .ZN(_01298_));
 NOR3_X4 _24256_ (.A1(_01140_),
    .A2(_01026_),
    .A3(_01225_),
    .ZN(_01299_));
 INV_X4 _24257_ (.A(_01059_),
    .ZN(_01300_));
 AOI21_X1 _24258_ (.A(_01143_),
    .B1(_01081_),
    .B2(_01300_),
    .ZN(_01301_));
 AOI21_X2 _24259_ (.A(_01299_),
    .B1(_01301_),
    .B2(_01116_),
    .ZN(_01302_));
 OAI221_X2 _24260_ (.A(_01240_),
    .B1(_01296_),
    .B2(_01298_),
    .C1(_01302_),
    .C2(_01184_),
    .ZN(_01303_));
 OAI22_X4 _24261_ (.A1(_01283_),
    .A2(_01276_),
    .B1(_01303_),
    .B2(_01294_),
    .ZN(_01304_));
 NOR2_X1 _24262_ (.A1(_15075_),
    .A2(_01006_),
    .ZN(_01305_));
 AOI21_X1 _24263_ (.A(_01305_),
    .B1(_01242_),
    .B2(_15078_),
    .ZN(_01306_));
 AOI21_X1 _24264_ (.A(_01096_),
    .B1(_01191_),
    .B2(_01306_),
    .ZN(_01307_));
 NOR3_X1 _24265_ (.A1(net923),
    .A2(_00979_),
    .A3(_01006_),
    .ZN(_01308_));
 NOR2_X4 _24266_ (.A1(_01084_),
    .A2(_01005_),
    .ZN(_01309_));
 AOI21_X4 _24267_ (.A(_01309_),
    .B1(_01005_),
    .B2(net8),
    .ZN(_01310_));
 NOR2_X1 _24268_ (.A1(net740),
    .A2(_01154_),
    .ZN(_01311_));
 AOI221_X2 _24269_ (.A(_01308_),
    .B1(_01310_),
    .B2(_01171_),
    .C1(net945),
    .C2(_01311_),
    .ZN(_01312_));
 OAI21_X2 _24270_ (.A(_01307_),
    .B1(_01191_),
    .B2(_01312_),
    .ZN(_01313_));
 OR2_X1 _24271_ (.A1(_01026_),
    .A2(_01139_),
    .ZN(_01314_));
 AND2_X1 _24272_ (.A1(_01201_),
    .A2(_01246_),
    .ZN(_01315_));
 OAI221_X2 _24273_ (.A(_01007_),
    .B1(_01223_),
    .B2(_01314_),
    .C1(_01315_),
    .C2(_00983_),
    .ZN(_01316_));
 NAND3_X1 _24274_ (.A1(net901),
    .A2(_01081_),
    .A3(_01160_),
    .ZN(_01317_));
 OR2_X1 _24275_ (.A1(_01212_),
    .A2(_01058_),
    .ZN(_01318_));
 MUX2_X1 _24276_ (.A(_00982_),
    .B(_01122_),
    .S(net844),
    .Z(_01319_));
 OAI221_X1 _24277_ (.A(_01317_),
    .B1(_01318_),
    .B2(_01172_),
    .C1(_01319_),
    .C2(_01118_),
    .ZN(_01320_));
 OAI21_X1 _24278_ (.A(_01316_),
    .B1(_01320_),
    .B2(_01007_),
    .ZN(_01321_));
 OAI21_X2 _24279_ (.A(_01313_),
    .B1(_01321_),
    .B2(_01151_),
    .ZN(_01322_));
 NAND2_X1 _24280_ (.A1(net923),
    .A2(_00978_),
    .ZN(_01323_));
 AND2_X1 _24281_ (.A1(_01080_),
    .A2(_01323_),
    .ZN(_01324_));
 AOI221_X2 _24282_ (.A(_01066_),
    .B1(_01231_),
    .B2(_01324_),
    .C1(_01146_),
    .C2(_15084_),
    .ZN(_01325_));
 AOI22_X1 _24283_ (.A1(_15073_),
    .A2(_01159_),
    .B1(_01083_),
    .B2(_01147_),
    .ZN(_01326_));
 NOR2_X1 _24284_ (.A1(_01096_),
    .A2(_01326_),
    .ZN(_01327_));
 OAI21_X1 _24285_ (.A(_01007_),
    .B1(_01325_),
    .B2(_01327_),
    .ZN(_01328_));
 AOI221_X1 _24286_ (.A(_01024_),
    .B1(_01105_),
    .B2(_01073_),
    .C1(_01315_),
    .C2(_01143_),
    .ZN(_01329_));
 NAND2_X1 _24287_ (.A1(_01159_),
    .A2(_01060_),
    .ZN(_01330_));
 OAI221_X1 _24288_ (.A(_01104_),
    .B1(_01107_),
    .B2(_01070_),
    .C1(_01330_),
    .C2(_00981_),
    .ZN(_01331_));
 AOI21_X1 _24289_ (.A(_01329_),
    .B1(_01331_),
    .B2(_01170_),
    .ZN(_01332_));
 OAI21_X1 _24290_ (.A(_01328_),
    .B1(_01332_),
    .B2(_01190_),
    .ZN(_01333_));
 AOI221_X2 _24291_ (.A(_01304_),
    .B1(_01322_),
    .B2(_01209_),
    .C1(_01219_),
    .C2(_01333_),
    .ZN(_00098_));
 NAND2_X1 _24292_ (.A1(_00988_),
    .A2(_01125_),
    .ZN(_01334_));
 NAND2_X1 _24293_ (.A1(_01172_),
    .A2(_01242_),
    .ZN(_01335_));
 OAI221_X1 _24294_ (.A(_01191_),
    .B1(_01310_),
    .B2(_01027_),
    .C1(_01335_),
    .C2(_01103_),
    .ZN(_01336_));
 OAI221_X1 _24295_ (.A(_01258_),
    .B1(_01335_),
    .B2(net682),
    .C1(_01300_),
    .C2(_00981_),
    .ZN(_01337_));
 AND3_X1 _24296_ (.A1(_01170_),
    .A2(_01336_),
    .A3(_01337_),
    .ZN(_01338_));
 AOI21_X1 _24297_ (.A(_01142_),
    .B1(_01164_),
    .B2(_01114_),
    .ZN(_01339_));
 AOI21_X2 _24298_ (.A(_01140_),
    .B1(_01060_),
    .B2(_01080_),
    .ZN(_01340_));
 AOI21_X1 _24299_ (.A(_01339_),
    .B1(_01340_),
    .B2(_00982_),
    .ZN(_01341_));
 NAND2_X1 _24300_ (.A1(net1056),
    .A2(_01107_),
    .ZN(_01342_));
 AOI21_X1 _24301_ (.A(_01242_),
    .B1(_01106_),
    .B2(_15061_),
    .ZN(_01343_));
 AOI221_X2 _24302_ (.A(_01096_),
    .B1(_01341_),
    .B2(_01242_),
    .C1(_01342_),
    .C2(_01343_),
    .ZN(_01344_));
 NAND4_X1 _24303_ (.A1(net844),
    .A2(_15050_),
    .A3(_01066_),
    .A4(_01091_),
    .ZN(_01345_));
 AOI22_X2 _24304_ (.A1(_00961_),
    .A2(_01142_),
    .B1(_01023_),
    .B2(net519),
    .ZN(_01346_));
 AOI21_X4 _24305_ (.A(_01091_),
    .B1(_01066_),
    .B2(_01118_),
    .ZN(_01347_));
 OAI221_X2 _24306_ (.A(_01345_),
    .B1(_01346_),
    .B2(_01122_),
    .C1(_01231_),
    .C2(_01347_),
    .ZN(_01348_));
 NAND2_X1 _24307_ (.A1(_01171_),
    .A2(_01023_),
    .ZN(_01349_));
 NAND2_X1 _24308_ (.A1(_01212_),
    .A2(_01066_),
    .ZN(_01350_));
 NAND2_X1 _24309_ (.A1(_01349_),
    .A2(_01350_),
    .ZN(_01351_));
 NOR3_X1 _24310_ (.A1(net741),
    .A2(_01143_),
    .A3(_01024_),
    .ZN(_01352_));
 AOI221_X2 _24311_ (.A(_01348_),
    .B1(_01351_),
    .B2(net743),
    .C1(_01258_),
    .C2(_01352_),
    .ZN(_01353_));
 OAI21_X1 _24312_ (.A(_01007_),
    .B1(_01160_),
    .B2(_01068_),
    .ZN(_01354_));
 OAI33_X1 _24313_ (.A1(_01344_),
    .A2(_01338_),
    .A3(_01334_),
    .B1(_01353_),
    .B2(_01354_),
    .B3(_01238_),
    .ZN(_01355_));
 NAND2_X1 _24314_ (.A1(_00988_),
    .A2(_01064_),
    .ZN(_01356_));
 NOR2_X4 _24315_ (.A1(_01241_),
    .A2(_01158_),
    .ZN(_01357_));
 NAND2_X2 _24316_ (.A1(_01066_),
    .A2(_01006_),
    .ZN(_01358_));
 NAND2_X2 _24317_ (.A1(_01087_),
    .A2(_00979_),
    .ZN(_01359_));
 OR2_X4 _24318_ (.A1(_01060_),
    .A2(_00979_),
    .ZN(_01360_));
 AOI21_X4 _24319_ (.A(_01099_),
    .B1(_01360_),
    .B2(_01359_),
    .ZN(_01361_));
 NOR3_X4 _24320_ (.A1(_01361_),
    .A2(_01358_),
    .A3(_01357_),
    .ZN(_01362_));
 NAND3_X1 _24321_ (.A1(net945),
    .A2(_01122_),
    .A3(_01154_),
    .ZN(_01363_));
 AOI21_X1 _24322_ (.A(_01067_),
    .B1(_01273_),
    .B2(_01363_),
    .ZN(_01364_));
 AOI21_X4 _24323_ (.A(_01309_),
    .B1(_01006_),
    .B2(_15050_),
    .ZN(_01365_));
 NAND2_X1 _24324_ (.A1(_01122_),
    .A2(_01154_),
    .ZN(_01366_));
 OAI221_X2 _24325_ (.A(_01143_),
    .B1(_01365_),
    .B2(_01158_),
    .C1(_01366_),
    .C2(net1056),
    .ZN(_01367_));
 OAI21_X1 _24326_ (.A(_15061_),
    .B1(_01027_),
    .B2(_01123_),
    .ZN(_01368_));
 AOI221_X2 _24327_ (.A(_01281_),
    .B1(_01082_),
    .B2(net740),
    .C1(_01108_),
    .C2(_01071_),
    .ZN(_01369_));
 AOI221_X2 _24328_ (.A(_01362_),
    .B1(_01367_),
    .B2(_01364_),
    .C1(_01368_),
    .C2(_01369_),
    .ZN(_01370_));
 NOR2_X2 _24329_ (.A1(_01370_),
    .A2(_01356_),
    .ZN(_01371_));
 NAND2_X1 _24330_ (.A1(_00989_),
    .A2(_01064_),
    .ZN(_01372_));
 OAI21_X1 _24331_ (.A(_01160_),
    .B1(net945),
    .B2(_01212_),
    .ZN(_01373_));
 AOI221_X2 _24332_ (.A(_01358_),
    .B1(_01373_),
    .B2(_01099_),
    .C1(_01105_),
    .C2(_01147_),
    .ZN(_01374_));
 AND2_X1 _24333_ (.A1(_01171_),
    .A2(_01114_),
    .ZN(_01375_));
 NOR2_X1 _24334_ (.A1(_00980_),
    .A2(_01140_),
    .ZN(_01376_));
 AOI221_X2 _24335_ (.A(_01293_),
    .B1(_01267_),
    .B2(_01375_),
    .C1(_01376_),
    .C2(_01274_),
    .ZN(_01377_));
 NAND3_X1 _24336_ (.A1(_01118_),
    .A2(_01052_),
    .A3(_01055_),
    .ZN(_01378_));
 AOI21_X1 _24337_ (.A(_01174_),
    .B1(_01378_),
    .B2(_01178_),
    .ZN(_01379_));
 NOR3_X1 _24338_ (.A1(_01027_),
    .A2(_01139_),
    .A3(_01175_),
    .ZN(_01380_));
 NAND2_X2 _24339_ (.A1(_01212_),
    .A2(_01225_),
    .ZN(_01381_));
 NAND2_X1 _24340_ (.A1(_01104_),
    .A2(_01381_),
    .ZN(_01382_));
 OAI33_X1 _24341_ (.A1(_01281_),
    .A2(_01379_),
    .A3(_01380_),
    .B1(_01299_),
    .B2(_01382_),
    .B3(_01184_),
    .ZN(_01383_));
 NOR4_X1 _24342_ (.A1(_01383_),
    .A2(_01374_),
    .A3(_01377_),
    .A4(_01372_),
    .ZN(_01384_));
 NAND2_X1 _24343_ (.A1(_01212_),
    .A2(_01091_),
    .ZN(_01385_));
 NOR2_X1 _24344_ (.A1(_00982_),
    .A2(_01197_),
    .ZN(_01386_));
 AOI21_X1 _24345_ (.A(_01119_),
    .B1(_01158_),
    .B2(_01211_),
    .ZN(_01387_));
 AOI221_X1 _24346_ (.A(_01024_),
    .B1(_01385_),
    .B2(_01386_),
    .C1(_01387_),
    .C2(_01174_),
    .ZN(_01388_));
 NAND3_X1 _24347_ (.A1(_01185_),
    .A2(_01201_),
    .A3(_01164_),
    .ZN(_01389_));
 OAI21_X1 _24348_ (.A(_01186_),
    .B1(_01258_),
    .B2(_01103_),
    .ZN(_01390_));
 OAI21_X1 _24349_ (.A(_01389_),
    .B1(_01390_),
    .B2(_01185_),
    .ZN(_01391_));
 AOI21_X1 _24350_ (.A(_01388_),
    .B1(_01391_),
    .B2(_01129_),
    .ZN(_01392_));
 NOR2_X1 _24351_ (.A1(_01220_),
    .A2(_01392_),
    .ZN(_01393_));
 NOR4_X2 _24352_ (.A1(_01384_),
    .A2(_01355_),
    .A3(_01371_),
    .A4(_01393_),
    .ZN(_00099_));
 NAND3_X1 _24353_ (.A1(_00981_),
    .A2(_01274_),
    .A3(_01246_),
    .ZN(_01394_));
 AND2_X1 _24354_ (.A1(_01067_),
    .A2(_01160_),
    .ZN(_01395_));
 NAND2_X1 _24355_ (.A1(_01027_),
    .A2(_01270_),
    .ZN(_01396_));
 OAI21_X1 _24356_ (.A(_01396_),
    .B1(_01258_),
    .B2(net925),
    .ZN(_01397_));
 AOI221_X1 _24357_ (.A(_01007_),
    .B1(_01394_),
    .B2(_01395_),
    .C1(_01397_),
    .C2(_01170_),
    .ZN(_01398_));
 AOI21_X1 _24358_ (.A(_00962_),
    .B1(_01026_),
    .B2(_01066_),
    .ZN(_01399_));
 OAI221_X2 _24359_ (.A(_01146_),
    .B1(_01399_),
    .B2(net901),
    .C1(_15050_),
    .C2(_01172_),
    .ZN(_01400_));
 NAND2_X1 _24360_ (.A1(net740),
    .A2(_01066_),
    .ZN(_01401_));
 OAI221_X2 _24361_ (.A(_01081_),
    .B1(_01349_),
    .B2(_01108_),
    .C1(_01401_),
    .C2(_01172_),
    .ZN(_01402_));
 MUX2_X1 _24362_ (.A(_01174_),
    .B(_01225_),
    .S(_01067_),
    .Z(_01403_));
 AOI221_X2 _24363_ (.A(_01156_),
    .B1(_01400_),
    .B2(_01402_),
    .C1(_01403_),
    .C2(net901),
    .ZN(_01404_));
 OAI21_X1 _24364_ (.A(_01209_),
    .B1(_01398_),
    .B2(_01404_),
    .ZN(_01405_));
 AOI21_X1 _24365_ (.A(_01026_),
    .B1(_01158_),
    .B2(_01047_),
    .ZN(_01406_));
 NAND2_X1 _24366_ (.A1(net836),
    .A2(_01081_),
    .ZN(_01407_));
 NOR2_X1 _24367_ (.A1(_00983_),
    .A2(net738),
    .ZN(_01408_));
 AOI221_X1 _24368_ (.A(_01096_),
    .B1(_01166_),
    .B2(_01406_),
    .C1(_01408_),
    .C2(_01407_),
    .ZN(_01409_));
 AOI21_X1 _24369_ (.A(net738),
    .B1(_01159_),
    .B2(_01147_),
    .ZN(_01410_));
 AOI221_X1 _24370_ (.A(_01068_),
    .B1(_01407_),
    .B2(_01273_),
    .C1(_01410_),
    .C2(_01144_),
    .ZN(_01411_));
 OAI21_X1 _24371_ (.A(_01190_),
    .B1(_01409_),
    .B2(_01411_),
    .ZN(_01412_));
 NOR2_X2 _24372_ (.A1(_15070_),
    .A2(_01228_),
    .ZN(_01413_));
 NOR2_X1 _24373_ (.A1(_01087_),
    .A2(_00979_),
    .ZN(_01414_));
 OR2_X1 _24374_ (.A1(_01068_),
    .A2(_01414_),
    .ZN(_01415_));
 OAI21_X1 _24375_ (.A(_01178_),
    .B1(_01258_),
    .B2(_01113_),
    .ZN(_01416_));
 OAI21_X1 _24376_ (.A(_01378_),
    .B1(_01091_),
    .B2(_01087_),
    .ZN(_01417_));
 MUX2_X1 _24377_ (.A(_01416_),
    .B(_01417_),
    .S(_01185_),
    .Z(_01418_));
 OAI221_X2 _24378_ (.A(_01156_),
    .B1(_01413_),
    .B2(_01415_),
    .C1(_01418_),
    .C2(_01129_),
    .ZN(_01419_));
 NAND3_X1 _24379_ (.A1(_01219_),
    .A2(_01412_),
    .A3(_01419_),
    .ZN(_01420_));
 NAND2_X1 _24380_ (.A1(_01125_),
    .A2(_01024_),
    .ZN(_01421_));
 NOR3_X1 _24381_ (.A1(_01212_),
    .A2(_01080_),
    .A3(_01154_),
    .ZN(_01422_));
 OAI21_X1 _24382_ (.A(_15050_),
    .B1(_00980_),
    .B2(_01422_),
    .ZN(_01423_));
 AOI21_X2 _24383_ (.A(_01005_),
    .B1(_01166_),
    .B2(net937),
    .ZN(_01424_));
 NOR2_X2 _24384_ (.A1(_01090_),
    .A2(_01153_),
    .ZN(_01425_));
 OAI21_X1 _24385_ (.A(net939),
    .B1(_01090_),
    .B2(_01005_),
    .ZN(_01426_));
 AOI221_X2 _24386_ (.A(_01424_),
    .B1(_01425_),
    .B2(_00961_),
    .C1(net8),
    .C2(_01426_),
    .ZN(_01427_));
 AOI221_X2 _24387_ (.A(_01421_),
    .B1(_01427_),
    .B2(_01423_),
    .C1(_01105_),
    .C2(net1056),
    .ZN(_01428_));
 MUX2_X1 _24388_ (.A(_01192_),
    .B(_01287_),
    .S(_01158_),
    .Z(_01429_));
 OAI21_X2 _24389_ (.A(_01025_),
    .B1(_01429_),
    .B2(_01007_),
    .ZN(_01430_));
 NOR3_X4 _24390_ (.A1(_01039_),
    .A2(_01300_),
    .A3(_01044_),
    .ZN(_01431_));
 NOR2_X2 _24391_ (.A1(_01431_),
    .A2(_01058_),
    .ZN(_01432_));
 OAI221_X2 _24392_ (.A(_01381_),
    .B1(_00981_),
    .B2(_01432_),
    .C1(_01092_),
    .C2(_01047_),
    .ZN(_01433_));
 AOI21_X2 _24393_ (.A(_01430_),
    .B1(_01190_),
    .B2(_01433_),
    .ZN(_01434_));
 OR3_X4 _24394_ (.A1(_01428_),
    .A2(_00989_),
    .A3(_01434_),
    .ZN(_01435_));
 AOI21_X1 _24395_ (.A(_01273_),
    .B1(_01106_),
    .B2(_15050_),
    .ZN(_01436_));
 OAI21_X1 _24396_ (.A(_01064_),
    .B1(_01358_),
    .B2(_01436_),
    .ZN(_01437_));
 NOR2_X1 _24397_ (.A1(_00982_),
    .A2(_01253_),
    .ZN(_01438_));
 NOR2_X2 _24398_ (.A1(_01142_),
    .A2(_01006_),
    .ZN(_01439_));
 NOR2_X1 _24399_ (.A1(_01431_),
    .A2(_01248_),
    .ZN(_01440_));
 OAI21_X1 _24400_ (.A(_01246_),
    .B1(_01099_),
    .B2(_01073_),
    .ZN(_01441_));
 AOI221_X2 _24401_ (.A(_01438_),
    .B1(_01439_),
    .B2(_01440_),
    .C1(_01174_),
    .C2(_01441_),
    .ZN(_01442_));
 AOI21_X1 _24402_ (.A(_01067_),
    .B1(_01440_),
    .B2(_01439_),
    .ZN(_01443_));
 NOR3_X2 _24403_ (.A1(_01143_),
    .A2(_01058_),
    .A3(_01140_),
    .ZN(_01444_));
 NOR3_X1 _24404_ (.A1(_01026_),
    .A2(_01075_),
    .A3(_01248_),
    .ZN(_01445_));
 NOR3_X1 _24405_ (.A1(_01096_),
    .A2(_01444_),
    .A3(_01445_),
    .ZN(_01446_));
 OR2_X1 _24406_ (.A1(_01443_),
    .A2(_01446_),
    .ZN(_01447_));
 AOI221_X2 _24407_ (.A(_01437_),
    .B1(_01442_),
    .B2(_01170_),
    .C1(_01447_),
    .C2(_01156_),
    .ZN(_01448_));
 OAI211_X2 _24408_ (.A(_01405_),
    .B(_01420_),
    .C1(_01448_),
    .C2(_01435_),
    .ZN(_00100_));
 OR2_X1 _24409_ (.A1(_01170_),
    .A2(_01098_),
    .ZN(_01449_));
 MUX2_X1 _24410_ (.A(_01211_),
    .B(_01074_),
    .S(_01174_),
    .Z(_01450_));
 OAI21_X1 _24411_ (.A(_01156_),
    .B1(_01450_),
    .B2(_01191_),
    .ZN(_01451_));
 AOI22_X1 _24412_ (.A1(net950),
    .A2(_01105_),
    .B1(_01417_),
    .B2(_01144_),
    .ZN(_01452_));
 OAI22_X1 _24413_ (.A1(_01449_),
    .A2(_01451_),
    .B1(_01452_),
    .B2(_01358_),
    .ZN(_01453_));
 OAI21_X1 _24414_ (.A(_01439_),
    .B1(_01197_),
    .B2(_01088_),
    .ZN(_01454_));
 OAI21_X1 _24415_ (.A(_01155_),
    .B1(_01146_),
    .B2(_01059_),
    .ZN(_01455_));
 AOI21_X1 _24416_ (.A(_01425_),
    .B1(_01455_),
    .B2(_01074_),
    .ZN(_01456_));
 AOI21_X1 _24417_ (.A(_01425_),
    .B1(_01106_),
    .B2(_01155_),
    .ZN(_01457_));
 OAI221_X2 _24418_ (.A(_01454_),
    .B1(_01456_),
    .B2(_15077_),
    .C1(_01284_),
    .C2(_01457_),
    .ZN(_01458_));
 NOR2_X1 _24419_ (.A1(_01151_),
    .A2(_01372_),
    .ZN(_01459_));
 AOI22_X1 _24420_ (.A1(_01209_),
    .A2(_01453_),
    .B1(_01458_),
    .B2(_01459_),
    .ZN(_01460_));
 MUX2_X1 _24421_ (.A(_01192_),
    .B(_01060_),
    .S(_01080_),
    .Z(_01461_));
 AOI221_X2 _24422_ (.A(_01242_),
    .B1(_01461_),
    .B2(_01143_),
    .C1(_01083_),
    .C2(_01147_),
    .ZN(_01462_));
 AOI221_X1 _24423_ (.A(_01155_),
    .B1(_01106_),
    .B2(_01192_),
    .C1(_01159_),
    .C2(_01103_),
    .ZN(_01463_));
 NOR3_X1 _24424_ (.A1(_01129_),
    .A2(_01462_),
    .A3(_01463_),
    .ZN(_01464_));
 AOI21_X1 _24425_ (.A(_01272_),
    .B1(_01122_),
    .B2(_01103_),
    .ZN(_01465_));
 NOR2_X1 _24426_ (.A1(_01119_),
    .A2(net737),
    .ZN(_01466_));
 MUX2_X1 _24427_ (.A(_01465_),
    .B(_01466_),
    .S(_00983_),
    .Z(_01467_));
 AOI21_X1 _24428_ (.A(_01159_),
    .B1(_00981_),
    .B2(_01073_),
    .ZN(_01468_));
 AOI21_X1 _24429_ (.A(_01468_),
    .B1(_01105_),
    .B2(_01211_),
    .ZN(_01469_));
 OAI22_X2 _24430_ (.A1(_01467_),
    .A2(_01293_),
    .B1(_01469_),
    .B2(_01184_),
    .ZN(_01470_));
 OAI21_X1 _24431_ (.A(_01240_),
    .B1(_01464_),
    .B2(_01470_),
    .ZN(_01471_));
 AOI21_X1 _24432_ (.A(_01144_),
    .B1(_01131_),
    .B2(_01163_),
    .ZN(_01472_));
 NOR2_X1 _24433_ (.A1(net741),
    .A2(_01261_),
    .ZN(_01473_));
 AOI21_X1 _24434_ (.A(_01144_),
    .B1(_01186_),
    .B2(_01202_),
    .ZN(_01474_));
 NOR2_X1 _24435_ (.A1(net682),
    .A2(_01109_),
    .ZN(_01475_));
 OAI33_X1 _24436_ (.A1(_01293_),
    .A2(_01472_),
    .A3(_01473_),
    .B1(_01474_),
    .B2(_01358_),
    .B3(_01475_),
    .ZN(_01476_));
 NAND2_X1 _24437_ (.A1(_01023_),
    .A2(_01080_),
    .ZN(_01477_));
 OAI221_X2 _24438_ (.A(_01155_),
    .B1(net686),
    .B2(_01477_),
    .C1(_01350_),
    .C2(_01092_),
    .ZN(_01478_));
 NAND2_X1 _24439_ (.A1(_01092_),
    .A2(_01401_),
    .ZN(_01479_));
 MUX2_X1 _24440_ (.A(_01158_),
    .B(_01196_),
    .S(_01023_),
    .Z(_01480_));
 AOI221_X2 _24441_ (.A(_01478_),
    .B1(_01479_),
    .B2(_15050_),
    .C1(net741),
    .C2(_01480_),
    .ZN(_01481_));
 OAI21_X1 _24442_ (.A(_01219_),
    .B1(_01481_),
    .B2(_01476_),
    .ZN(_01482_));
 XNOR2_X1 _24443_ (.A(_15061_),
    .B(_01242_),
    .ZN(_01483_));
 AOI22_X2 _24444_ (.A1(_01074_),
    .A2(_01083_),
    .B1(_01071_),
    .B2(_01192_),
    .ZN(_01484_));
 OAI221_X2 _24445_ (.A(_01151_),
    .B1(_01261_),
    .B2(_01483_),
    .C1(_01484_),
    .C2(_01156_),
    .ZN(_01485_));
 NAND2_X1 _24446_ (.A1(_01155_),
    .A2(_01116_),
    .ZN(_01486_));
 AOI21_X1 _24447_ (.A(net950),
    .B1(_01210_),
    .B2(_01486_),
    .ZN(_01487_));
 OAI21_X1 _24448_ (.A(_01267_),
    .B1(_01091_),
    .B2(net924),
    .ZN(_01488_));
 NOR2_X2 _24449_ (.A1(_01026_),
    .A2(net737),
    .ZN(_01489_));
 AOI221_X1 _24450_ (.A(_01242_),
    .B1(_01488_),
    .B2(_01026_),
    .C1(_01489_),
    .C2(_01385_),
    .ZN(_01490_));
 AOI221_X1 _24451_ (.A(_01154_),
    .B1(_01106_),
    .B2(_01070_),
    .C1(_01465_),
    .C2(_00980_),
    .ZN(_01491_));
 OR2_X1 _24452_ (.A1(_01490_),
    .A2(_01491_),
    .ZN(_01492_));
 OAI221_X2 _24453_ (.A(_01183_),
    .B1(_01485_),
    .B2(_01487_),
    .C1(_01492_),
    .C2(_01151_),
    .ZN(_01493_));
 AND4_X2 _24454_ (.A1(_01460_),
    .A2(_01471_),
    .A3(_01482_),
    .A4(_01493_),
    .ZN(_00101_));
 INV_X2 _24455_ (.A(_01087_),
    .ZN(_01494_));
 MUX2_X1 _24456_ (.A(_01494_),
    .B(_01103_),
    .S(_01099_),
    .Z(_01495_));
 AOI221_X2 _24457_ (.A(_01068_),
    .B1(_01071_),
    .B2(net901),
    .C1(_01495_),
    .C2(_01185_),
    .ZN(_01496_));
 NAND2_X1 _24458_ (.A1(_01190_),
    .A2(_01286_),
    .ZN(_01497_));
 OAI21_X1 _24459_ (.A(_01129_),
    .B1(_01475_),
    .B2(_01339_),
    .ZN(_01498_));
 AOI21_X1 _24460_ (.A(_01170_),
    .B1(_01258_),
    .B2(_15072_),
    .ZN(_01499_));
 OAI21_X1 _24461_ (.A(_01359_),
    .B1(_15077_),
    .B2(net901),
    .ZN(_01500_));
 OAI21_X1 _24462_ (.A(_01499_),
    .B1(_01500_),
    .B2(_01258_),
    .ZN(_01501_));
 NAND2_X1 _24463_ (.A1(_01498_),
    .A2(_01501_),
    .ZN(_01502_));
 OAI221_X2 _24464_ (.A(_01240_),
    .B1(_01496_),
    .B2(_01497_),
    .C1(_01502_),
    .C2(_01190_),
    .ZN(_01503_));
 OR3_X1 _24465_ (.A1(_15071_),
    .A2(_15080_),
    .A3(_01122_),
    .ZN(_01504_));
 MUX2_X1 _24466_ (.A(_00962_),
    .B(_00982_),
    .S(_01212_),
    .Z(_01505_));
 OAI21_X1 _24467_ (.A(_01504_),
    .B1(_01505_),
    .B2(_01146_),
    .ZN(_01506_));
 AND2_X1 _24468_ (.A1(_01297_),
    .A2(_01506_),
    .ZN(_01507_));
 OAI21_X1 _24469_ (.A(_01270_),
    .B1(_01122_),
    .B2(_01047_),
    .ZN(_01508_));
 AOI221_X1 _24470_ (.A(_01184_),
    .B1(_01508_),
    .B2(_01143_),
    .C1(_01105_),
    .C2(net925),
    .ZN(_01509_));
 MUX2_X1 _24471_ (.A(_01211_),
    .B(_01494_),
    .S(_00979_),
    .Z(_01510_));
 OAI21_X2 _24472_ (.A(_01266_),
    .B1(_01081_),
    .B2(_01510_),
    .ZN(_01511_));
 AOI221_X2 _24473_ (.A(_01097_),
    .B1(_01055_),
    .B2(_01052_),
    .C1(_01192_),
    .C2(_01026_),
    .ZN(_01512_));
 OAI21_X1 _24474_ (.A(_01270_),
    .B1(_01158_),
    .B2(net945),
    .ZN(_01513_));
 OAI21_X1 _24475_ (.A(_01378_),
    .B1(_01060_),
    .B2(_01099_),
    .ZN(_01514_));
 MUX2_X1 _24476_ (.A(_01513_),
    .B(_01514_),
    .S(_00980_),
    .Z(_01515_));
 OAI22_X2 _24477_ (.A1(_01511_),
    .A2(_01512_),
    .B1(_01515_),
    .B2(_01293_),
    .ZN(_01516_));
 OR4_X4 _24478_ (.A1(_01372_),
    .A2(_01516_),
    .A3(_01509_),
    .A4(_01507_),
    .ZN(_01517_));
 OAI21_X1 _24479_ (.A(_01323_),
    .B1(_00981_),
    .B2(_01084_),
    .ZN(_01518_));
 MUX2_X1 _24480_ (.A(_15073_),
    .B(_01518_),
    .S(_01191_),
    .Z(_01519_));
 OAI21_X1 _24481_ (.A(_15070_),
    .B1(_01140_),
    .B2(_01213_),
    .ZN(_01520_));
 AOI21_X1 _24482_ (.A(_01281_),
    .B1(_01148_),
    .B2(_15077_),
    .ZN(_01521_));
 AOI22_X2 _24483_ (.A1(_01245_),
    .A2(_01519_),
    .B1(_01520_),
    .B2(_01521_),
    .ZN(_01522_));
 NOR3_X1 _24484_ (.A1(_15077_),
    .A2(_01222_),
    .A3(_01061_),
    .ZN(_01523_));
 NOR3_X1 _24485_ (.A1(_15070_),
    .A2(_01140_),
    .A3(_01225_),
    .ZN(_01524_));
 OAI21_X1 _24486_ (.A(_01266_),
    .B1(_01523_),
    .B2(_01524_),
    .ZN(_01525_));
 MUX2_X1 _24487_ (.A(_01103_),
    .B(net741),
    .S(_01159_),
    .Z(_01526_));
 OAI221_X1 _24488_ (.A(_01252_),
    .B1(_01526_),
    .B2(_15070_),
    .C1(_01109_),
    .C2(_01147_),
    .ZN(_01527_));
 NAND4_X2 _24489_ (.A1(_01219_),
    .A2(_01522_),
    .A3(_01525_),
    .A4(_01527_),
    .ZN(_01528_));
 AOI22_X1 _24490_ (.A1(_01147_),
    .A2(_01083_),
    .B1(_01071_),
    .B2(net950),
    .ZN(_01529_));
 OAI21_X1 _24491_ (.A(net741),
    .B1(_15070_),
    .B2(_01225_),
    .ZN(_01530_));
 NAND3_X1 _24492_ (.A1(_01151_),
    .A2(_01529_),
    .A3(_01530_),
    .ZN(_01531_));
 AOI22_X1 _24493_ (.A1(net950),
    .A2(_01185_),
    .B1(_01106_),
    .B2(_01211_),
    .ZN(_01532_));
 NAND3_X1 _24494_ (.A1(_01129_),
    .A2(_01381_),
    .A3(_01532_),
    .ZN(_01533_));
 AOI21_X1 _24495_ (.A(_01190_),
    .B1(_01531_),
    .B2(_01533_),
    .ZN(_01534_));
 OR2_X1 _24496_ (.A1(_01172_),
    .A2(_01417_),
    .ZN(_01535_));
 AOI21_X1 _24497_ (.A(_01024_),
    .B1(_01105_),
    .B2(_15050_),
    .ZN(_01536_));
 NAND2_X1 _24498_ (.A1(_01284_),
    .A2(_00980_),
    .ZN(_01537_));
 NAND3_X1 _24499_ (.A1(_01146_),
    .A2(_01160_),
    .A3(_01537_),
    .ZN(_01538_));
 OAI21_X1 _24500_ (.A(_01538_),
    .B1(_01191_),
    .B2(_01233_),
    .ZN(_01539_));
 AOI221_X2 _24501_ (.A(_01155_),
    .B1(_01535_),
    .B2(_01536_),
    .C1(_01539_),
    .C2(_01170_),
    .ZN(_01540_));
 OAI21_X2 _24502_ (.A(_01183_),
    .B1(_01540_),
    .B2(_01534_),
    .ZN(_01541_));
 NAND4_X4 _24503_ (.A1(_01503_),
    .A2(_01517_),
    .A3(_01528_),
    .A4(_01541_),
    .ZN(_00102_));
 NOR2_X2 _24504_ (.A1(net739),
    .A2(_01156_),
    .ZN(_01542_));
 OAI21_X2 _24505_ (.A(_01542_),
    .B1(_01505_),
    .B2(_01191_),
    .ZN(_01543_));
 OAI21_X1 _24506_ (.A(_01270_),
    .B1(_01159_),
    .B2(_01192_),
    .ZN(_01544_));
 OAI21_X1 _24507_ (.A(_01144_),
    .B1(_01191_),
    .B2(_01060_),
    .ZN(_01545_));
 OAI221_X2 _24508_ (.A(_01156_),
    .B1(_01544_),
    .B2(_01144_),
    .C1(_01545_),
    .C2(_01123_),
    .ZN(_01546_));
 AOI21_X2 _24509_ (.A(_01151_),
    .B1(_01543_),
    .B2(_01546_),
    .ZN(_01547_));
 OAI21_X1 _24510_ (.A(_01027_),
    .B1(_01139_),
    .B2(_01175_),
    .ZN(_01548_));
 AND3_X1 _24511_ (.A1(_01155_),
    .A2(_01257_),
    .A3(_01548_),
    .ZN(_01549_));
 AOI21_X1 _24512_ (.A(_01142_),
    .B1(_01091_),
    .B2(_01300_),
    .ZN(_01550_));
 AOI221_X2 _24513_ (.A(_01154_),
    .B1(_01274_),
    .B2(_01550_),
    .C1(_01174_),
    .C2(_01108_),
    .ZN(_01551_));
 NOR3_X2 _24514_ (.A1(_01549_),
    .A2(_01129_),
    .A3(_01551_),
    .ZN(_01552_));
 NOR3_X1 _24515_ (.A1(_01372_),
    .A2(_01547_),
    .A3(_01552_),
    .ZN(_01553_));
 AOI21_X1 _24516_ (.A(_01083_),
    .B1(_01258_),
    .B2(_01068_),
    .ZN(_01554_));
 OAI22_X1 _24517_ (.A1(_15070_),
    .A2(_01170_),
    .B1(_01554_),
    .B2(_01070_),
    .ZN(_01555_));
 AOI22_X4 _24518_ (.A1(_01018_),
    .A2(_01021_),
    .B1(_01052_),
    .B2(_01055_),
    .ZN(_01556_));
 AOI21_X1 _24519_ (.A(_01119_),
    .B1(_01556_),
    .B2(_01147_),
    .ZN(_01557_));
 NOR2_X1 _24520_ (.A1(_15077_),
    .A2(_01557_),
    .ZN(_01558_));
 OAI21_X1 _24521_ (.A(_01190_),
    .B1(_01555_),
    .B2(_01558_),
    .ZN(_01559_));
 NOR2_X1 _24522_ (.A1(_00962_),
    .A2(_01171_),
    .ZN(_01560_));
 NOR2_X1 _24523_ (.A1(_01192_),
    .A2(_01143_),
    .ZN(_01561_));
 NOR2_X1 _24524_ (.A1(_01023_),
    .A2(_01122_),
    .ZN(_01562_));
 AOI221_X2 _24525_ (.A(_01242_),
    .B1(_01560_),
    .B2(_01556_),
    .C1(_01561_),
    .C2(_01562_),
    .ZN(_01563_));
 NOR3_X1 _24526_ (.A1(net742),
    .A2(_01024_),
    .A3(_01146_),
    .ZN(_01564_));
 AOI21_X1 _24527_ (.A(_01564_),
    .B1(_01191_),
    .B2(_01096_),
    .ZN(_01565_));
 AOI21_X1 _24528_ (.A(_01105_),
    .B1(_01562_),
    .B2(_15070_),
    .ZN(_01566_));
 OAI221_X2 _24529_ (.A(_01563_),
    .B1(_01565_),
    .B2(_15050_),
    .C1(net901),
    .C2(_01566_),
    .ZN(_01567_));
 AOI21_X1 _24530_ (.A(_01334_),
    .B1(_01559_),
    .B2(_01567_),
    .ZN(_01568_));
 OAI222_X2 _24531_ (.A1(net950),
    .A2(_01092_),
    .B1(_01109_),
    .B2(_01113_),
    .C1(_01084_),
    .C2(_01107_),
    .ZN(_01569_));
 OAI21_X1 _24532_ (.A(_01185_),
    .B1(_01196_),
    .B2(_01248_),
    .ZN(_01570_));
 AOI21_X1 _24533_ (.A(_01184_),
    .B1(_01406_),
    .B2(_01166_),
    .ZN(_01571_));
 AOI22_X1 _24534_ (.A1(_01252_),
    .A2(_01569_),
    .B1(_01570_),
    .B2(_01571_),
    .ZN(_01572_));
 OAI21_X1 _24535_ (.A(_01160_),
    .B1(_01144_),
    .B2(net901),
    .ZN(_01573_));
 AOI21_X1 _24536_ (.A(_01511_),
    .B1(_01573_),
    .B2(_01258_),
    .ZN(_01574_));
 AOI21_X1 _24537_ (.A(_01272_),
    .B1(_01159_),
    .B2(net901),
    .ZN(_01575_));
 OAI22_X1 _24538_ (.A1(net1056),
    .A2(_01210_),
    .B1(_01575_),
    .B2(_01185_),
    .ZN(_01576_));
 AOI21_X1 _24539_ (.A(_01574_),
    .B1(_01576_),
    .B2(_01297_),
    .ZN(_01577_));
 AOI21_X1 _24540_ (.A(_01356_),
    .B1(_01572_),
    .B2(_01577_),
    .ZN(_01578_));
 NOR2_X1 _24541_ (.A1(_01067_),
    .A2(_01188_),
    .ZN(_01579_));
 NOR2_X1 _24542_ (.A1(net737),
    .A2(_01223_),
    .ZN(_01580_));
 OAI21_X2 _24543_ (.A(_01579_),
    .B1(_01580_),
    .B2(_01027_),
    .ZN(_01581_));
 OAI21_X1 _24544_ (.A(_01091_),
    .B1(_01287_),
    .B2(_01414_),
    .ZN(_01582_));
 OAI21_X1 _24545_ (.A(_01582_),
    .B1(_01099_),
    .B2(_15080_),
    .ZN(_01583_));
 AOI21_X1 _24546_ (.A(_01155_),
    .B1(_01583_),
    .B2(_01067_),
    .ZN(_01584_));
 AOI21_X1 _24547_ (.A(_01197_),
    .B1(_01099_),
    .B2(_01147_),
    .ZN(_01585_));
 OAI21_X1 _24548_ (.A(_01024_),
    .B1(_01585_),
    .B2(_01172_),
    .ZN(_01586_));
 AOI21_X1 _24549_ (.A(_01248_),
    .B1(_01083_),
    .B2(net925),
    .ZN(_01587_));
 OAI22_X1 _24550_ (.A1(_01438_),
    .A2(_01586_),
    .B1(_01587_),
    .B2(_01096_),
    .ZN(_01588_));
 AOI221_X1 _24551_ (.A(_01238_),
    .B1(_01581_),
    .B2(_01584_),
    .C1(_01588_),
    .C2(_01156_),
    .ZN(_01589_));
 NOR4_X1 _24552_ (.A1(_01578_),
    .A2(_01568_),
    .A3(_01553_),
    .A4(_01589_),
    .ZN(_00103_));
 INV_X1 _24553_ (.A(_06466_),
    .ZN(_01590_));
 NOR2_X1 _24554_ (.A1(_01590_),
    .A2(_08975_),
    .ZN(_01591_));
 NOR2_X1 _24555_ (.A1(_06466_),
    .A2(_08975_),
    .ZN(_01592_));
 XOR2_X2 _24556_ (.A(\sa30_sub[1] ),
    .B(\sa01_sr[1] ),
    .Z(_01593_));
 XNOR2_X2 _24557_ (.A(_09796_),
    .B(_09799_),
    .ZN(_01594_));
 XNOR2_X2 _24558_ (.A(_01594_),
    .B(_01593_),
    .ZN(_01595_));
 XOR2_X1 _24559_ (.A(\sa30_sub[0] ),
    .B(\sa21_sr[0] ),
    .Z(_01596_));
 XNOR2_X1 _24560_ (.A(_01596_),
    .B(\sa11_sr[1] ),
    .ZN(_01597_));
 XNOR2_X2 _24561_ (.A(_01597_),
    .B(_01595_),
    .ZN(_01598_));
 MUX2_X2 _24562_ (.A(_01591_),
    .B(_01592_),
    .S(_01598_),
    .Z(_01599_));
 NAND3_X1 _24563_ (.A1(_06466_),
    .A2(_09180_),
    .A3(_00467_),
    .ZN(_01600_));
 NAND2_X2 _24564_ (.A1(_01590_),
    .A2(_09818_),
    .ZN(_01601_));
 OAI21_X4 _24565_ (.A(_01600_),
    .B1(_00467_),
    .B2(_01601_),
    .ZN(_01602_));
 NOR2_X4 _24566_ (.A1(_01602_),
    .A2(_01599_),
    .ZN(_01603_));
 INV_X8 _24567_ (.A(_01603_),
    .ZN(_01604_));
 BUF_X4 clone254 (.A(net807),
    .Z(net806));
 BUF_X32 _24569_ (.A(_01604_),
    .Z(_15092_));
 XNOR2_X1 _24570_ (.A(\sa11_sr[0] ),
    .B(_01594_),
    .ZN(_01606_));
 NAND3_X1 _24571_ (.A1(_06451_),
    .A2(_09118_),
    .A3(_12517_),
    .ZN(_01607_));
 NOR2_X1 _24572_ (.A1(_06451_),
    .A2(_08994_),
    .ZN(_01608_));
 NAND2_X1 _24573_ (.A1(_12510_),
    .A2(_01608_),
    .ZN(_01609_));
 AOI21_X1 _24574_ (.A(_01606_),
    .B1(_01607_),
    .B2(_01609_),
    .ZN(_01610_));
 XOR2_X1 _24575_ (.A(\sa11_sr[0] ),
    .B(_01594_),
    .Z(_01611_));
 NAND2_X1 _24576_ (.A1(_12517_),
    .A2(_01608_),
    .ZN(_01612_));
 NAND3_X1 _24577_ (.A1(_06451_),
    .A2(_09116_),
    .A3(_12510_),
    .ZN(_01613_));
 AOI21_X1 _24578_ (.A(_01611_),
    .B1(_01612_),
    .B2(_01613_),
    .ZN(_01614_));
 INV_X1 _24579_ (.A(_06451_),
    .ZN(_01615_));
 NAND3_X1 _24580_ (.A1(_01615_),
    .A2(_09179_),
    .A3(_00468_),
    .ZN(_01616_));
 NAND2_X1 _24581_ (.A1(_06451_),
    .A2(_09103_),
    .ZN(_01617_));
 OAI21_X1 _24582_ (.A(_01616_),
    .B1(_01617_),
    .B2(_00468_),
    .ZN(_01618_));
 OR3_X4 _24583_ (.A1(_01610_),
    .A2(_01614_),
    .A3(_01618_),
    .ZN(_01619_));
 INV_X4 _24584_ (.A(_01619_),
    .ZN(_15097_));
 XOR2_X2 _24585_ (.A(net636),
    .B(_09762_),
    .Z(_01620_));
 XOR2_X1 _24586_ (.A(\sa30_sub[1] ),
    .B(_01620_),
    .Z(_01621_));
 NAND3_X1 _24587_ (.A1(_06483_),
    .A2(_09195_),
    .A3(_12535_),
    .ZN(_01622_));
 NOR2_X1 _24588_ (.A1(_06483_),
    .A2(_09727_),
    .ZN(_01623_));
 NAND2_X1 _24589_ (.A1(_12529_),
    .A2(_01623_),
    .ZN(_01624_));
 AOI21_X2 _24590_ (.A(_01621_),
    .B1(_01622_),
    .B2(_01624_),
    .ZN(_01625_));
 XNOR2_X1 _24591_ (.A(net755),
    .B(_01620_),
    .ZN(_01626_));
 NAND2_X1 _24592_ (.A1(_12535_),
    .A2(_01623_),
    .ZN(_01627_));
 NAND3_X1 _24593_ (.A1(_06483_),
    .A2(_09856_),
    .A3(_12529_),
    .ZN(_01628_));
 AOI21_X2 _24594_ (.A(_01626_),
    .B1(_01627_),
    .B2(_01628_),
    .ZN(_01629_));
 NAND3_X1 _24595_ (.A1(_06486_),
    .A2(_11938_),
    .A3(_00469_),
    .ZN(_01630_));
 NAND2_X1 _24596_ (.A1(_06483_),
    .A2(_11938_),
    .ZN(_01631_));
 OAI21_X2 _24597_ (.A(_01630_),
    .B1(_01631_),
    .B2(_00469_),
    .ZN(_01632_));
 NOR3_X4 _24598_ (.A1(_01625_),
    .A2(_01629_),
    .A3(_01632_),
    .ZN(_01633_));
 INV_X1 _24599_ (.A(_01633_),
    .ZN(_01634_));
 BUF_X4 _24600_ (.A(_01634_),
    .Z(_01635_));
 BUF_X4 _24601_ (.A(_01635_),
    .Z(_01636_));
 BUF_X4 _24602_ (.A(_01636_),
    .Z(_01637_));
 BUF_X4 _24603_ (.A(_01637_),
    .Z(_15113_));
 BUF_X8 _24604_ (.A(_01603_),
    .Z(_15087_));
 BUF_X4 _24605_ (.A(_01633_),
    .Z(_01638_));
 BUF_X4 _24606_ (.A(_01638_),
    .Z(_01639_));
 BUF_X4 _24607_ (.A(_01639_),
    .Z(_01640_));
 BUF_X4 _24608_ (.A(_01640_),
    .Z(_15106_));
 NAND2_X1 _24609_ (.A1(_06543_),
    .A2(_09158_),
    .ZN(_01641_));
 INV_X1 _24610_ (.A(_06543_),
    .ZN(_01642_));
 NAND2_X1 _24611_ (.A1(_01642_),
    .A2(_09158_),
    .ZN(_01643_));
 XNOR2_X1 _24612_ (.A(_09872_),
    .B(_09785_),
    .ZN(_01644_));
 XNOR2_X2 _24613_ (.A(_12615_),
    .B(_01644_),
    .ZN(_01645_));
 MUX2_X2 _24614_ (.A(_01641_),
    .B(_01643_),
    .S(_01645_),
    .Z(_01646_));
 NOR3_X2 _24615_ (.A1(_01642_),
    .A2(_09158_),
    .A3(\text_in_r[77] ),
    .ZN(_01647_));
 NOR2_X1 _24616_ (.A1(_06543_),
    .A2(_09803_),
    .ZN(_01648_));
 AOI21_X4 _24617_ (.A(_01647_),
    .B1(_01648_),
    .B2(\text_in_r[77] ),
    .ZN(_01649_));
 AND2_X1 _24618_ (.A1(_01646_),
    .A2(_01649_),
    .ZN(_01650_));
 BUF_X4 _24619_ (.A(_01650_),
    .Z(_01651_));
 BUF_X4 _24620_ (.A(_01651_),
    .Z(_01652_));
 XNOR2_X1 _24621_ (.A(_09809_),
    .B(_09786_),
    .ZN(_01653_));
 XNOR2_X2 _24622_ (.A(_12629_),
    .B(_01653_),
    .ZN(_01654_));
 MUX2_X2 _24623_ (.A(\text_in_r[78] ),
    .B(_01654_),
    .S(_09803_),
    .Z(_01655_));
 XOR2_X2 _24624_ (.A(_06556_),
    .B(_01655_),
    .Z(_01656_));
 XNOR2_X1 _24625_ (.A(_09787_),
    .B(_09799_),
    .ZN(_01657_));
 XNOR2_X2 _24626_ (.A(_09790_),
    .B(_09742_),
    .ZN(_01658_));
 XNOR2_X1 _24627_ (.A(_01657_),
    .B(_01658_),
    .ZN(_01659_));
 MUX2_X2 _24628_ (.A(\text_in_r[79] ),
    .B(_01659_),
    .S(_09158_),
    .Z(_01660_));
 XNOR2_X2 _24629_ (.A(_06565_),
    .B(_01660_),
    .ZN(_01661_));
 NOR2_X2 _24630_ (.A1(_01656_),
    .A2(_01661_),
    .ZN(_01662_));
 NAND2_X1 _24631_ (.A1(_01652_),
    .A2(_01662_),
    .ZN(_01663_));
 INV_X1 _24632_ (.A(_06528_),
    .ZN(_01664_));
 NOR2_X1 _24633_ (.A1(net951),
    .A2(\text_in_r[76] ),
    .ZN(_01665_));
 XNOR2_X1 _24634_ (.A(_09813_),
    .B(_09799_),
    .ZN(_01666_));
 XNOR2_X1 _24635_ (.A(_09841_),
    .B(_09808_),
    .ZN(_01667_));
 XNOR2_X2 _24636_ (.A(_01666_),
    .B(_01667_),
    .ZN(_01668_));
 XOR2_X2 _24637_ (.A(_12557_),
    .B(_01668_),
    .Z(_01669_));
 AOI211_X2 _24638_ (.A(_01664_),
    .B(_01665_),
    .C1(_01669_),
    .C2(_09175_),
    .ZN(_01670_));
 NAND2_X2 _24639_ (.A1(_08974_),
    .A2(\text_in_r[76] ),
    .ZN(_01671_));
 INV_X1 _24640_ (.A(_01671_),
    .ZN(_01672_));
 XNOR2_X2 _24641_ (.A(_12557_),
    .B(_01668_),
    .ZN(_01673_));
 AOI211_X2 _24642_ (.A(_06528_),
    .B(_01672_),
    .C1(_01673_),
    .C2(_09175_),
    .ZN(_01674_));
 NAND2_X1 _24643_ (.A1(_06511_),
    .A2(_09175_),
    .ZN(_01675_));
 INV_X1 _24644_ (.A(_06511_),
    .ZN(_01676_));
 NAND2_X1 _24645_ (.A1(_01676_),
    .A2(_09138_),
    .ZN(_01677_));
 XNOR2_X1 _24646_ (.A(_09868_),
    .B(_09799_),
    .ZN(_01678_));
 XNOR2_X1 _24647_ (.A(_09759_),
    .B(_09839_),
    .ZN(_01679_));
 XNOR2_X2 _24648_ (.A(_01678_),
    .B(_01679_),
    .ZN(_01680_));
 XNOR2_X1 _24649_ (.A(_09763_),
    .B(_12575_),
    .ZN(_01681_));
 XNOR2_X2 _24650_ (.A(_01680_),
    .B(_01681_),
    .ZN(_01682_));
 MUX2_X1 _24651_ (.A(_01675_),
    .B(_01677_),
    .S(_01682_),
    .Z(_01683_));
 BUF_X8 _24652_ (.A(_01683_),
    .Z(_01684_));
 BUF_X8 _24653_ (.A(_01684_),
    .Z(_01685_));
 OR3_X2 _24654_ (.A1(_01676_),
    .A2(_09116_),
    .A3(\text_in_r[75] ),
    .ZN(_01686_));
 NAND3_X2 _24655_ (.A1(_01676_),
    .A2(_09180_),
    .A3(\text_in_r[75] ),
    .ZN(_01687_));
 AND2_X1 _24656_ (.A1(_01686_),
    .A2(_01687_),
    .ZN(_01688_));
 BUF_X8 _24657_ (.A(_01688_),
    .Z(_01689_));
 BUF_X8 _24658_ (.A(_01689_),
    .Z(_01690_));
 AOI211_X2 _24659_ (.A(_01670_),
    .B(_01674_),
    .C1(_01685_),
    .C2(_01690_),
    .ZN(_01691_));
 AOI21_X1 _24660_ (.A(_01663_),
    .B1(_01691_),
    .B2(_15111_),
    .ZN(_01692_));
 NOR2_X1 _24661_ (.A1(_01676_),
    .A2(_08995_),
    .ZN(_01693_));
 NOR2_X1 _24662_ (.A1(_06511_),
    .A2(_08995_),
    .ZN(_01694_));
 MUX2_X1 _24663_ (.A(_01693_),
    .B(_01694_),
    .S(_01682_),
    .Z(_01695_));
 BUF_X4 _24664_ (.A(_01695_),
    .Z(_01696_));
 NAND2_X4 _24665_ (.A1(_01686_),
    .A2(_01687_),
    .ZN(_01697_));
 NOR2_X2 _24666_ (.A1(_01696_),
    .A2(_01697_),
    .ZN(_01698_));
 BUF_X4 _24667_ (.A(_01698_),
    .Z(_01699_));
 BUF_X4 _24668_ (.A(_01699_),
    .Z(_01700_));
 BUF_X4 _24669_ (.A(_01700_),
    .Z(_01701_));
 NOR2_X1 _24670_ (.A1(_01670_),
    .A2(_01674_),
    .ZN(_01702_));
 BUF_X4 _24671_ (.A(_01702_),
    .Z(_01703_));
 BUF_X4 _24672_ (.A(_01703_),
    .Z(_01704_));
 BUF_X4 _24673_ (.A(_01704_),
    .Z(_01705_));
 BUF_X4 _24674_ (.A(_15089_),
    .Z(_01706_));
 INV_X8 _24675_ (.A(_01706_),
    .ZN(_01707_));
 NOR2_X4 _24676_ (.A1(_01633_),
    .A2(_01707_),
    .ZN(_01708_));
 NAND2_X1 _24677_ (.A1(_01705_),
    .A2(net757),
    .ZN(_01709_));
 OR2_X1 _24678_ (.A1(_09803_),
    .A2(\text_in_r[76] ),
    .ZN(_01710_));
 OAI211_X4 _24679_ (.A(_06528_),
    .B(_01710_),
    .C1(_01673_),
    .C2(_09136_),
    .ZN(_01711_));
 OAI211_X4 _24680_ (.A(_01664_),
    .B(_01671_),
    .C1(_01669_),
    .C2(_09136_),
    .ZN(_01712_));
 NAND2_X4 _24681_ (.A1(_01711_),
    .A2(_01712_),
    .ZN(_01713_));
 INV_X2 _24682_ (.A(_15093_),
    .ZN(_01714_));
 MUX2_X2 _24683_ (.A(_15095_),
    .B(_01714_),
    .S(_01638_),
    .Z(_01715_));
 NAND2_X1 _24684_ (.A1(_01713_),
    .A2(_01715_),
    .ZN(_01716_));
 NAND2_X1 _24685_ (.A1(_01709_),
    .A2(_01716_),
    .ZN(_01717_));
 BUF_X4 _24686_ (.A(_15088_),
    .Z(_01718_));
 BUF_X4 _24687_ (.A(_01696_),
    .Z(_01719_));
 BUF_X4 _24688_ (.A(_01697_),
    .Z(_01720_));
 OAI21_X2 _24689_ (.A(_01638_),
    .B1(_01719_),
    .B2(_01720_),
    .ZN(_01721_));
 CLKBUF_X3 _24690_ (.A(_01721_),
    .Z(_01722_));
 AOI21_X4 _24691_ (.A(_01619_),
    .B1(_01684_),
    .B2(_01689_),
    .ZN(_01723_));
 BUF_X4 _24692_ (.A(_01699_),
    .Z(_01724_));
 CLKBUF_X3 _24693_ (.A(_15090_),
    .Z(_01725_));
 AOI21_X1 _24694_ (.A(_01723_),
    .B1(_01724_),
    .B2(_01725_),
    .ZN(_01726_));
 OAI22_X1 _24695_ (.A1(_01718_),
    .A2(_01722_),
    .B1(_01726_),
    .B2(_15106_),
    .ZN(_01727_));
 BUF_X4 _24696_ (.A(_01713_),
    .Z(_01728_));
 CLKBUF_X3 _24697_ (.A(_01728_),
    .Z(_01729_));
 AOI22_X1 _24698_ (.A1(_01701_),
    .A2(_01717_),
    .B1(_01727_),
    .B2(_01729_),
    .ZN(_01730_));
 NAND2_X1 _24699_ (.A1(_01692_),
    .A2(_01730_),
    .ZN(_01731_));
 BUF_X4 _24700_ (.A(_01652_),
    .Z(_01732_));
 XNOR2_X2 _24701_ (.A(_06556_),
    .B(_01655_),
    .ZN(_01733_));
 BUF_X4 _24702_ (.A(_01733_),
    .Z(_01734_));
 BUF_X4 _24703_ (.A(_01734_),
    .Z(_01735_));
 XOR2_X2 _24704_ (.A(_06565_),
    .B(_01660_),
    .Z(_01736_));
 NAND2_X1 _24705_ (.A1(_01735_),
    .A2(_01736_),
    .ZN(_01737_));
 NOR2_X1 _24706_ (.A1(_01732_),
    .A2(_01737_),
    .ZN(_01738_));
 BUF_X4 _24707_ (.A(_01703_),
    .Z(_01739_));
 BUF_X4 _24708_ (.A(_01739_),
    .Z(_01740_));
 AOI21_X4 _24709_ (.A(net1127),
    .B1(_01684_),
    .B2(_01689_),
    .ZN(_01741_));
 AOI21_X2 _24710_ (.A(_01741_),
    .B1(_01699_),
    .B2(_01725_),
    .ZN(_01742_));
 BUF_X4 _24711_ (.A(_01635_),
    .Z(_01743_));
 NAND2_X4 _24712_ (.A1(_01684_),
    .A2(_01689_),
    .ZN(_01744_));
 NAND2_X2 _24713_ (.A1(_01743_),
    .A2(_01744_),
    .ZN(_01745_));
 BUF_X2 _24714_ (.A(_15100_),
    .Z(_01746_));
 INV_X2 _24715_ (.A(_01746_),
    .ZN(_01747_));
 OAI22_X2 _24716_ (.A1(_15113_),
    .A2(_01742_),
    .B1(_01745_),
    .B2(_01747_),
    .ZN(_01748_));
 NOR2_X1 _24717_ (.A1(_01740_),
    .A2(_01748_),
    .ZN(_01749_));
 BUF_X4 _24718_ (.A(_01638_),
    .Z(_01750_));
 BUF_X4 _24719_ (.A(_15093_),
    .Z(_01751_));
 NAND3_X2 _24720_ (.A1(_01751_),
    .A2(_01685_),
    .A3(_01690_),
    .ZN(_01752_));
 INV_X2 _24721_ (.A(_01725_),
    .ZN(_01753_));
 BUF_X4 _24722_ (.A(_01696_),
    .Z(_01754_));
 BUF_X4 _24723_ (.A(_01697_),
    .Z(_01755_));
 OAI21_X1 _24724_ (.A(_01753_),
    .B1(_01754_),
    .B2(_01755_),
    .ZN(_01756_));
 AND3_X2 _24725_ (.A1(_01750_),
    .A2(_01752_),
    .A3(_01756_),
    .ZN(_01757_));
 NAND3_X4 _24726_ (.A1(_01635_),
    .A2(_01685_),
    .A3(_01690_),
    .ZN(_01758_));
 BUF_X4 _24727_ (.A(_15098_),
    .Z(_01759_));
 OAI21_X1 _24728_ (.A(_01705_),
    .B1(_01758_),
    .B2(net1133),
    .ZN(_01760_));
 NOR2_X1 _24729_ (.A1(_01757_),
    .A2(_01760_),
    .ZN(_01761_));
 OAI21_X1 _24730_ (.A(_01738_),
    .B1(_01749_),
    .B2(_01761_),
    .ZN(_01762_));
 NAND2_X2 _24731_ (.A1(_01646_),
    .A2(_01649_),
    .ZN(_01763_));
 NAND2_X2 _24732_ (.A1(_01763_),
    .A2(_01713_),
    .ZN(_01764_));
 NAND2_X2 _24733_ (.A1(_01718_),
    .A2(_01743_),
    .ZN(_01765_));
 NAND2_X1 _24734_ (.A1(net1133),
    .A2(_01640_),
    .ZN(_01766_));
 AOI21_X1 _24735_ (.A(_01724_),
    .B1(_01765_),
    .B2(_01766_),
    .ZN(_01767_));
 BUF_X4 _24736_ (.A(_01744_),
    .Z(_01768_));
 BUF_X4 _24737_ (.A(_01768_),
    .Z(_01769_));
 BUF_X4 clone126 (.A(_01603_),
    .Z(net126));
 BUF_X4 _24739_ (.A(_15102_),
    .Z(_01771_));
 BUF_X4 _24740_ (.A(_01743_),
    .Z(_01772_));
 NAND2_X1 _24741_ (.A1(_01771_),
    .A2(_01772_),
    .ZN(_01773_));
 BUF_X16 _24742_ (.A(_01707_),
    .Z(_01774_));
 NAND2_X1 _24743_ (.A1(_01774_),
    .A2(_01640_),
    .ZN(_01775_));
 AOI21_X1 _24744_ (.A(_01769_),
    .B1(_01773_),
    .B2(_01775_),
    .ZN(_01776_));
 NOR3_X1 _24745_ (.A1(_01764_),
    .A2(_01767_),
    .A3(_01776_),
    .ZN(_01777_));
 NAND2_X1 _24746_ (.A1(_01734_),
    .A2(_01661_),
    .ZN(_01778_));
 NOR2_X1 _24747_ (.A1(_01777_),
    .A2(_01778_),
    .ZN(_01779_));
 OAI22_X1 _24748_ (.A1(_01774_),
    .A2(_01721_),
    .B1(_01758_),
    .B2(_01759_),
    .ZN(_01780_));
 AOI21_X4 _24749_ (.A(_01633_),
    .B1(_01684_),
    .B2(_01689_),
    .ZN(_01781_));
 NOR3_X4 _24750_ (.A1(_01634_),
    .A2(_01696_),
    .A3(_01697_),
    .ZN(_01782_));
 OR2_X2 _24751_ (.A1(_01781_),
    .A2(_01782_),
    .ZN(_01783_));
 INV_X1 _24752_ (.A(_01718_),
    .ZN(_01784_));
 AOI21_X1 _24753_ (.A(_01780_),
    .B1(_01783_),
    .B2(_01784_),
    .ZN(_01785_));
 NAND3_X4 _24754_ (.A1(_01706_),
    .A2(_01684_),
    .A3(_01689_),
    .ZN(_01786_));
 BUF_X4 _24755_ (.A(_01743_),
    .Z(_01787_));
 AOI21_X2 _24756_ (.A(_01786_),
    .B1(_01787_),
    .B2(net125),
    .ZN(_01788_));
 BUF_X8 _24757_ (.A(_01706_),
    .Z(_01789_));
 NOR2_X2 _24758_ (.A1(net806),
    .A2(_01750_),
    .ZN(_01790_));
 BUF_X4 _24759_ (.A(_01603_),
    .Z(_01791_));
 BUF_X4 _24760_ (.A(_01698_),
    .Z(_01792_));
 BUF_X4 _24761_ (.A(_01792_),
    .Z(_01793_));
 NAND2_X1 _24762_ (.A1(_01791_),
    .A2(_01793_),
    .ZN(_01794_));
 AOI21_X1 _24763_ (.A(_01788_),
    .B1(_01790_),
    .B2(_01794_),
    .ZN(_01795_));
 MUX2_X1 _24764_ (.A(_01785_),
    .B(_01795_),
    .S(_01739_),
    .Z(_01796_));
 BUF_X4 _24765_ (.A(_01763_),
    .Z(_01797_));
 BUF_X4 _24766_ (.A(_01797_),
    .Z(_01798_));
 BUF_X4 _24767_ (.A(_01763_),
    .Z(_01799_));
 NAND2_X2 _24768_ (.A1(_01799_),
    .A2(_01704_),
    .ZN(_01800_));
 CLKBUF_X3 _24769_ (.A(_01769_),
    .Z(_01801_));
 BUF_X8 _24770_ (.A(_01619_),
    .Z(_01802_));
 NOR2_X4 _24771_ (.A1(_01802_),
    .A2(_01635_),
    .ZN(_01803_));
 AOI21_X2 _24772_ (.A(_01803_),
    .B1(_01802_),
    .B2(net125),
    .ZN(_01804_));
 XNOR2_X1 _24773_ (.A(_01801_),
    .B(_01804_),
    .ZN(_01805_));
 OAI221_X1 _24774_ (.A(_01779_),
    .B1(_01796_),
    .B2(_01798_),
    .C1(_01800_),
    .C2(_01805_),
    .ZN(_01806_));
 BUF_X4 _24775_ (.A(_01656_),
    .Z(_01807_));
 BUF_X4 _24776_ (.A(_01736_),
    .Z(_01808_));
 BUF_X4 _24777_ (.A(_01746_),
    .Z(_01809_));
 NAND4_X1 _24778_ (.A1(_01809_),
    .A2(_01640_),
    .A3(_01793_),
    .A4(_01704_),
    .ZN(_01810_));
 MUX2_X1 _24779_ (.A(_01774_),
    .B(_01771_),
    .S(_01713_),
    .Z(_01811_));
 OAI21_X2 _24780_ (.A(_01810_),
    .B1(_01811_),
    .B2(_01722_),
    .ZN(_01812_));
 OAI21_X4 _24781_ (.A(_01802_),
    .B1(_01754_),
    .B2(_01755_),
    .ZN(_01813_));
 NOR2_X1 _24782_ (.A1(_01704_),
    .A2(_01813_),
    .ZN(_01814_));
 INV_X8 _24783_ (.A(net756),
    .ZN(_01815_));
 NAND3_X4 _24784_ (.A1(_01815_),
    .A2(_01685_),
    .A3(_01690_),
    .ZN(_01816_));
 NAND2_X1 _24785_ (.A1(_01772_),
    .A2(_01816_),
    .ZN(_01817_));
 OAI21_X1 _24786_ (.A(_01652_),
    .B1(_01814_),
    .B2(_01817_),
    .ZN(_01818_));
 AOI211_X2 _24787_ (.A(_01743_),
    .B(_01723_),
    .C1(_01699_),
    .C2(net125),
    .ZN(_01819_));
 OAI21_X2 _24788_ (.A(_01759_),
    .B1(_01719_),
    .B2(_01720_),
    .ZN(_01820_));
 AOI21_X1 _24789_ (.A(_01640_),
    .B1(_01786_),
    .B2(_01820_),
    .ZN(_01821_));
 NOR3_X1 _24790_ (.A1(_01739_),
    .A2(_01819_),
    .A3(_01821_),
    .ZN(_01822_));
 BUF_X4 _24791_ (.A(_01768_),
    .Z(_01823_));
 NAND2_X2 _24792_ (.A1(_01753_),
    .A2(_01639_),
    .ZN(_01824_));
 AOI21_X1 _24793_ (.A(_01823_),
    .B1(_01765_),
    .B2(_01824_),
    .ZN(_01825_));
 BUF_X8 _24794_ (.A(_15095_),
    .Z(_01826_));
 OAI21_X1 _24795_ (.A(_01704_),
    .B1(_01722_),
    .B2(_01826_),
    .ZN(_01827_));
 OAI21_X1 _24796_ (.A(_01797_),
    .B1(_01825_),
    .B2(_01827_),
    .ZN(_01828_));
 OAI221_X2 _24797_ (.A(_01808_),
    .B1(_01812_),
    .B2(_01818_),
    .C1(_01822_),
    .C2(_01828_),
    .ZN(_01829_));
 BUF_X4 _24798_ (.A(_01728_),
    .Z(_01830_));
 OAI21_X1 _24799_ (.A(_01787_),
    .B1(_01602_),
    .B2(net593),
    .ZN(_01831_));
 NAND3_X1 _24800_ (.A1(_01724_),
    .A2(_01824_),
    .A3(_01831_),
    .ZN(_01832_));
 NOR2_X1 _24801_ (.A1(_01802_),
    .A2(_01639_),
    .ZN(_01833_));
 NOR2_X1 _24802_ (.A1(_01771_),
    .A2(_01787_),
    .ZN(_01834_));
 OAI21_X1 _24803_ (.A(_01769_),
    .B1(_01833_),
    .B2(_01834_),
    .ZN(_01835_));
 NAND4_X1 _24804_ (.A1(_01652_),
    .A2(_01830_),
    .A3(_01832_),
    .A4(_01835_),
    .ZN(_01836_));
 NOR2_X2 _24805_ (.A1(_01651_),
    .A2(_01713_),
    .ZN(_01837_));
 BUF_X4 _24806_ (.A(_01639_),
    .Z(_01838_));
 NAND3_X4 _24807_ (.A1(_01802_),
    .A2(_01685_),
    .A3(_01690_),
    .ZN(_01839_));
 OAI21_X4 _24808_ (.A(_01774_),
    .B1(_01719_),
    .B2(_01720_),
    .ZN(_01840_));
 NAND3_X1 _24809_ (.A1(_01838_),
    .A2(_01839_),
    .A3(_01840_),
    .ZN(_01841_));
 BUF_X4 _24810_ (.A(_01787_),
    .Z(_01842_));
 BUF_X2 clone162 (.A(net509),
    .Z(net162));
 INV_X4 _24812_ (.A(_15104_),
    .ZN(_01844_));
 OAI21_X1 _24813_ (.A(_01844_),
    .B1(_01754_),
    .B2(_01755_),
    .ZN(_01845_));
 NAND3_X1 _24814_ (.A1(_01842_),
    .A2(_01752_),
    .A3(_01845_),
    .ZN(_01846_));
 NAND3_X1 _24815_ (.A1(_01837_),
    .A2(_01841_),
    .A3(_01846_),
    .ZN(_01847_));
 NOR2_X1 _24816_ (.A1(_01652_),
    .A2(_01739_),
    .ZN(_01848_));
 NOR2_X1 _24817_ (.A1(net761),
    .A2(_01722_),
    .ZN(_01849_));
 OAI21_X2 _24818_ (.A(_01751_),
    .B1(_01719_),
    .B2(_01720_),
    .ZN(_01850_));
 AOI21_X1 _24819_ (.A(_01838_),
    .B1(_01839_),
    .B2(_01850_),
    .ZN(_01851_));
 OAI21_X1 _24820_ (.A(_01848_),
    .B1(_01849_),
    .B2(_01851_),
    .ZN(_01852_));
 NAND4_X4 _24821_ (.A1(_01646_),
    .A2(_01649_),
    .A3(_01711_),
    .A4(_01712_),
    .ZN(_01853_));
 NOR3_X4 _24822_ (.A1(_01751_),
    .A2(_01719_),
    .A3(_01720_),
    .ZN(_01854_));
 NOR4_X1 _24823_ (.A1(_01640_),
    .A2(_01723_),
    .A3(_01853_),
    .A4(_01854_),
    .ZN(_01855_));
 NOR2_X1 _24824_ (.A1(_01842_),
    .A2(_01853_),
    .ZN(_01856_));
 MUX2_X1 _24825_ (.A(_01844_),
    .B(_01791_),
    .S(_01699_),
    .Z(_01857_));
 AOI21_X1 _24826_ (.A(_01855_),
    .B1(_01856_),
    .B2(_01857_),
    .ZN(_01858_));
 NAND4_X2 _24827_ (.A1(_01836_),
    .A2(_01847_),
    .A3(_01852_),
    .A4(_01858_),
    .ZN(_01859_));
 OAI211_X2 _24828_ (.A(_01807_),
    .B(_01829_),
    .C1(_01859_),
    .C2(_01808_),
    .ZN(_01860_));
 AND4_X2 _24829_ (.A1(_01806_),
    .A2(_01762_),
    .A3(_01731_),
    .A4(_01860_),
    .ZN(_00104_));
 BUF_X8 _24830_ (.A(_01802_),
    .Z(_15086_));
 NOR2_X2 _24831_ (.A1(_01734_),
    .A2(_01661_),
    .ZN(_01861_));
 AOI21_X4 _24832_ (.A(_01706_),
    .B1(_01684_),
    .B2(_01689_),
    .ZN(_01862_));
 AOI21_X1 _24833_ (.A(_01862_),
    .B1(_01699_),
    .B2(_01826_),
    .ZN(_01863_));
 OAI221_X1 _24834_ (.A(_01799_),
    .B1(_01745_),
    .B2(_01771_),
    .C1(_01863_),
    .C2(_01772_),
    .ZN(_01864_));
 OAI21_X2 _24835_ (.A(_15097_),
    .B1(_01719_),
    .B2(_01720_),
    .ZN(_01865_));
 OAI22_X1 _24836_ (.A1(_01604_),
    .A2(_01865_),
    .B1(_01758_),
    .B2(_01774_),
    .ZN(_01866_));
 AOI21_X1 _24837_ (.A(_01866_),
    .B1(_01783_),
    .B2(_15086_),
    .ZN(_01867_));
 OAI221_X1 _24838_ (.A(_01864_),
    .B1(_01674_),
    .B2(_01670_),
    .C1(_01797_),
    .C2(_01867_),
    .ZN(_01868_));
 NOR3_X4 _24839_ (.A1(_01718_),
    .A2(_01696_),
    .A3(_01697_),
    .ZN(_01869_));
 OAI21_X1 _24840_ (.A(_01750_),
    .B1(_01862_),
    .B2(_01869_),
    .ZN(_01870_));
 NOR3_X2 _24841_ (.A1(_01802_),
    .A2(_01754_),
    .A3(_01755_),
    .ZN(_01871_));
 AOI21_X4 _24842_ (.A(_01815_),
    .B1(_01684_),
    .B2(_01689_),
    .ZN(_01872_));
 OAI21_X1 _24843_ (.A(_01787_),
    .B1(_01871_),
    .B2(net805),
    .ZN(_01873_));
 NAND3_X1 _24844_ (.A1(_01651_),
    .A2(_01870_),
    .A3(_01873_),
    .ZN(_01874_));
 MUX2_X1 _24845_ (.A(_01771_),
    .B(net125),
    .S(_01744_),
    .Z(_01875_));
 OAI221_X1 _24846_ (.A(_01799_),
    .B1(_01745_),
    .B2(_01844_),
    .C1(_01875_),
    .C2(_01772_),
    .ZN(_01876_));
 NAND3_X1 _24847_ (.A1(_01739_),
    .A2(_01874_),
    .A3(_01876_),
    .ZN(_01877_));
 AND3_X1 _24848_ (.A1(_01861_),
    .A2(_01868_),
    .A3(_01877_),
    .ZN(_01878_));
 NOR2_X1 _24849_ (.A1(_01826_),
    .A2(_01638_),
    .ZN(_01879_));
 INV_X1 _24850_ (.A(_01602_),
    .ZN(_01880_));
 NAND2_X1 _24851_ (.A1(_06466_),
    .A2(_11207_),
    .ZN(_01881_));
 NAND2_X1 _24852_ (.A1(_01590_),
    .A2(_11207_),
    .ZN(_01882_));
 MUX2_X2 _24853_ (.A(_01881_),
    .B(_01882_),
    .S(_01598_),
    .Z(_01883_));
 AOI21_X4 _24854_ (.A(_01635_),
    .B1(_01880_),
    .B2(_01883_),
    .ZN(_01884_));
 OR3_X1 _24855_ (.A1(_01713_),
    .A2(_01879_),
    .A3(_01884_),
    .ZN(_01885_));
 AOI21_X2 _24856_ (.A(_01768_),
    .B1(_01885_),
    .B2(_01716_),
    .ZN(_01886_));
 NAND2_X1 _24857_ (.A1(_15104_),
    .A2(_01638_),
    .ZN(_01887_));
 NOR2_X2 _24858_ (.A1(_01702_),
    .A2(_01708_),
    .ZN(_01888_));
 AOI221_X2 _24859_ (.A(_01698_),
    .B1(_01888_),
    .B2(_01887_),
    .C1(_01703_),
    .C2(_15118_),
    .ZN(_01889_));
 OR3_X4 _24860_ (.A1(_01889_),
    .A2(_01886_),
    .A3(_01797_),
    .ZN(_01890_));
 NAND3_X1 _24861_ (.A1(_01838_),
    .A2(_01816_),
    .A3(_01840_),
    .ZN(_01891_));
 NOR3_X4 _24862_ (.A1(_15097_),
    .A2(_01696_),
    .A3(_01697_),
    .ZN(_01892_));
 OAI21_X1 _24863_ (.A(_01637_),
    .B1(_01723_),
    .B2(_01892_),
    .ZN(_01893_));
 NAND2_X1 _24864_ (.A1(_01891_),
    .A2(_01893_),
    .ZN(_01894_));
 NAND2_X2 _24865_ (.A1(_15097_),
    .A2(_01793_),
    .ZN(_01895_));
 AOI21_X1 _24866_ (.A(_01741_),
    .B1(_01700_),
    .B2(_15092_),
    .ZN(_01896_));
 BUF_X4 _24867_ (.A(_01750_),
    .Z(_01897_));
 OAI22_X2 _24868_ (.A1(_15092_),
    .A2(_01895_),
    .B1(_01896_),
    .B2(_01897_),
    .ZN(_01898_));
 OAI221_X2 _24869_ (.A(_01890_),
    .B1(_01894_),
    .B2(_01800_),
    .C1(_01898_),
    .C2(_01764_),
    .ZN(_01899_));
 INV_X2 _24870_ (.A(_15102_),
    .ZN(_01900_));
 NOR3_X4 _24871_ (.A1(_01900_),
    .A2(_01696_),
    .A3(_01697_),
    .ZN(_01901_));
 OAI21_X1 _24872_ (.A(_01638_),
    .B1(net1132),
    .B2(_01901_),
    .ZN(_01902_));
 AOI21_X1 _24873_ (.A(_01763_),
    .B1(_01892_),
    .B2(_01635_),
    .ZN(_01903_));
 NOR3_X4 _24874_ (.A1(_01872_),
    .A2(_01892_),
    .A3(_01635_),
    .ZN(_01904_));
 AOI21_X1 _24875_ (.A(_01869_),
    .B1(_01744_),
    .B2(_01604_),
    .ZN(_01905_));
 AOI21_X2 _24876_ (.A(_01904_),
    .B1(_01905_),
    .B2(_01743_),
    .ZN(_01906_));
 AOI221_X2 _24877_ (.A(_01703_),
    .B1(_01902_),
    .B2(_01903_),
    .C1(_01906_),
    .C2(_01799_),
    .ZN(_01907_));
 NAND3_X2 _24878_ (.A1(_01636_),
    .A2(_01839_),
    .A3(_01840_),
    .ZN(_01908_));
 NAND3_X2 _24879_ (.A1(_01753_),
    .A2(_01685_),
    .A3(_01690_),
    .ZN(_01909_));
 OAI21_X1 _24880_ (.A(_01909_),
    .B1(_01699_),
    .B2(_01784_),
    .ZN(_01910_));
 OAI21_X1 _24881_ (.A(_01908_),
    .B1(_01910_),
    .B2(_01772_),
    .ZN(_01911_));
 NOR3_X2 _24882_ (.A1(_01844_),
    .A2(_01719_),
    .A3(_01720_),
    .ZN(_01912_));
 NOR3_X1 _24883_ (.A1(_01636_),
    .A2(net1130),
    .A3(_01912_),
    .ZN(_01913_));
 OAI21_X2 _24884_ (.A(_15102_),
    .B1(_01719_),
    .B2(_01720_),
    .ZN(_01914_));
 NAND2_X1 _24885_ (.A1(_01909_),
    .A2(_01914_),
    .ZN(_01915_));
 AOI21_X1 _24886_ (.A(_01913_),
    .B1(_01915_),
    .B2(_01772_),
    .ZN(_01916_));
 OAI22_X1 _24887_ (.A1(_01800_),
    .A2(_01911_),
    .B1(_01916_),
    .B2(_01853_),
    .ZN(_01917_));
 OR3_X2 _24888_ (.A1(_01735_),
    .A2(_01907_),
    .A3(_01917_),
    .ZN(_01918_));
 OAI21_X1 _24889_ (.A(_01772_),
    .B1(_01741_),
    .B2(_01869_),
    .ZN(_01919_));
 NAND3_X1 _24890_ (.A1(_01750_),
    .A2(_01839_),
    .A3(_01914_),
    .ZN(_01920_));
 AND3_X1 _24891_ (.A1(_01837_),
    .A2(_01919_),
    .A3(_01920_),
    .ZN(_01921_));
 MUX2_X1 _24892_ (.A(_01759_),
    .B(_15102_),
    .S(_01638_),
    .Z(_01922_));
 NOR2_X2 _24893_ (.A1(_01922_),
    .A2(_01768_),
    .ZN(_01923_));
 NOR3_X1 _24894_ (.A1(_15114_),
    .A2(_01799_),
    .A3(_01793_),
    .ZN(_01924_));
 NOR3_X1 _24895_ (.A1(_01739_),
    .A2(_01923_),
    .A3(_01924_),
    .ZN(_01925_));
 NOR2_X2 _24896_ (.A1(_01763_),
    .A2(_01713_),
    .ZN(_01926_));
 XNOR2_X2 _24897_ (.A(_01604_),
    .B(_01792_),
    .ZN(_01927_));
 AND3_X1 _24898_ (.A1(_01637_),
    .A2(_01926_),
    .A3(_01927_),
    .ZN(_01928_));
 NOR3_X1 _24899_ (.A1(_01921_),
    .A2(_01925_),
    .A3(_01928_),
    .ZN(_01929_));
 NOR2_X1 _24900_ (.A1(_01892_),
    .A2(_01872_),
    .ZN(_01930_));
 AOI21_X1 _24901_ (.A(_01807_),
    .B1(_01856_),
    .B2(_01930_),
    .ZN(_01931_));
 AOI21_X1 _24902_ (.A(_01808_),
    .B1(_01929_),
    .B2(_01931_),
    .ZN(_01932_));
 AOI221_X2 _24903_ (.A(_01878_),
    .B1(_01899_),
    .B2(_01662_),
    .C1(_01918_),
    .C2(_01932_),
    .ZN(_00105_));
 NAND3_X1 _24904_ (.A1(_01791_),
    .A2(_01802_),
    .A3(_01651_),
    .ZN(_01933_));
 NAND2_X1 _24905_ (.A1(_01823_),
    .A2(_01933_),
    .ZN(_01934_));
 MUX2_X1 _24906_ (.A(_01751_),
    .B(net763),
    .S(_01651_),
    .Z(_01935_));
 AOI221_X2 _24907_ (.A(_01934_),
    .B1(_01935_),
    .B2(_01838_),
    .C1(_01797_),
    .C2(_01790_),
    .ZN(_01936_));
 NOR2_X1 _24908_ (.A1(_15114_),
    .A2(_01797_),
    .ZN(_01937_));
 AOI21_X1 _24909_ (.A(_01937_),
    .B1(_01798_),
    .B2(_15111_),
    .ZN(_01938_));
 OAI21_X1 _24910_ (.A(_01729_),
    .B1(_01938_),
    .B2(_01801_),
    .ZN(_01939_));
 AOI21_X2 _24911_ (.A(_01862_),
    .B1(_01699_),
    .B2(_01718_),
    .ZN(_01940_));
 INV_X4 _24912_ (.A(_01759_),
    .ZN(_01941_));
 MUX2_X1 _24913_ (.A(_01941_),
    .B(net763),
    .S(_01792_),
    .Z(_01942_));
 MUX2_X1 _24914_ (.A(_01940_),
    .B(_01942_),
    .S(_01838_),
    .Z(_01943_));
 NOR3_X1 _24915_ (.A1(_01604_),
    .A2(_01792_),
    .A3(_01803_),
    .ZN(_01944_));
 MUX2_X1 _24916_ (.A(_01635_),
    .B(_01792_),
    .S(_01604_),
    .Z(_01945_));
 AOI221_X2 _24917_ (.A(_01944_),
    .B1(_01884_),
    .B2(_01865_),
    .C1(_01789_),
    .C2(_01945_),
    .ZN(_01946_));
 MUX2_X1 _24918_ (.A(_01943_),
    .B(_01946_),
    .S(_01798_),
    .Z(_01947_));
 OAI221_X2 _24919_ (.A(_01861_),
    .B1(_01936_),
    .B2(_01939_),
    .C1(_01947_),
    .C2(_01729_),
    .ZN(_01948_));
 OAI21_X1 _24920_ (.A(_01839_),
    .B1(_01700_),
    .B2(_01809_),
    .ZN(_01949_));
 NAND3_X4 _24921_ (.A1(_01844_),
    .A2(_01685_),
    .A3(_01690_),
    .ZN(_01950_));
 OAI21_X1 _24922_ (.A(_01950_),
    .B1(_01700_),
    .B2(_01791_),
    .ZN(_01951_));
 MUX2_X1 _24923_ (.A(_01949_),
    .B(_01951_),
    .S(_01842_),
    .Z(_01952_));
 OAI21_X1 _24924_ (.A(_01950_),
    .B1(_01700_),
    .B2(_01826_),
    .ZN(_01953_));
 OAI21_X1 _24925_ (.A(_01813_),
    .B1(_01823_),
    .B2(_01809_),
    .ZN(_01954_));
 MUX2_X1 _24926_ (.A(_01953_),
    .B(_01954_),
    .S(_01838_),
    .Z(_01955_));
 AOI22_X1 _24927_ (.A1(_01837_),
    .A2(_01952_),
    .B1(_01955_),
    .B2(_01926_),
    .ZN(_01956_));
 NAND3_X2 _24928_ (.A1(_01746_),
    .A2(_01684_),
    .A3(_01689_),
    .ZN(_01957_));
 AND2_X1 _24929_ (.A1(_01840_),
    .A2(_01957_),
    .ZN(_01958_));
 OAI21_X1 _24930_ (.A(_01841_),
    .B1(_01958_),
    .B2(_01897_),
    .ZN(_01959_));
 AOI21_X4 _24931_ (.A(_01743_),
    .B1(_01744_),
    .B2(_01604_),
    .ZN(_01960_));
 AOI21_X1 _24932_ (.A(_01879_),
    .B1(_01957_),
    .B2(_01960_),
    .ZN(_01961_));
 MUX2_X1 _24933_ (.A(_01959_),
    .B(_01961_),
    .S(_01652_),
    .Z(_01962_));
 OAI21_X2 _24934_ (.A(_01956_),
    .B1(_01962_),
    .B2(_01740_),
    .ZN(_01963_));
 NAND2_X1 _24935_ (.A1(_01807_),
    .A2(_01661_),
    .ZN(_01964_));
 BUF_X4 _24936_ (.A(_01661_),
    .Z(_01965_));
 NAND2_X1 _24937_ (.A1(_01604_),
    .A2(_01639_),
    .ZN(_01966_));
 OAI221_X2 _24938_ (.A(_01966_),
    .B1(_01755_),
    .B2(_01754_),
    .C1(_01714_),
    .C2(_01750_),
    .ZN(_01967_));
 AOI21_X1 _24939_ (.A(_01799_),
    .B1(_01793_),
    .B2(_15120_),
    .ZN(_01968_));
 NOR3_X4 _24940_ (.A1(_01638_),
    .A2(_01719_),
    .A3(_01720_),
    .ZN(_01969_));
 NAND2_X4 _24941_ (.A1(_01753_),
    .A2(_01815_),
    .ZN(_01970_));
 AOI21_X4 _24942_ (.A(_01970_),
    .B1(_01690_),
    .B2(_01685_),
    .ZN(_01971_));
 AOI22_X2 _24943_ (.A1(net1133),
    .A2(_01969_),
    .B1(_01971_),
    .B2(_01639_),
    .ZN(_01972_));
 NOR2_X1 _24944_ (.A1(_01781_),
    .A2(_01782_),
    .ZN(_01973_));
 OAI21_X2 _24945_ (.A(_01972_),
    .B1(_01973_),
    .B2(_01900_),
    .ZN(_01974_));
 AOI221_X2 _24946_ (.A(_01830_),
    .B1(_01967_),
    .B2(_01968_),
    .C1(_01974_),
    .C2(_01797_),
    .ZN(_01975_));
 AOI221_X2 _24947_ (.A(_01651_),
    .B1(_01781_),
    .B2(net761),
    .C1(_01940_),
    .C2(_01640_),
    .ZN(_01976_));
 BUF_X4 _24948_ (.A(_01768_),
    .Z(_01977_));
 NAND2_X1 _24949_ (.A1(_15109_),
    .A2(_01977_),
    .ZN(_01978_));
 NAND2_X1 _24950_ (.A1(_01751_),
    .A2(_01969_),
    .ZN(_01979_));
 AOI21_X1 _24951_ (.A(_01798_),
    .B1(_01978_),
    .B2(_01979_),
    .ZN(_01980_));
 NOR3_X1 _24952_ (.A1(_01740_),
    .A2(_01976_),
    .A3(_01980_),
    .ZN(_01981_));
 NOR3_X2 _24953_ (.A1(_01975_),
    .A2(_01965_),
    .A3(_01981_),
    .ZN(_01982_));
 AOI21_X1 _24954_ (.A(_01637_),
    .B1(_01865_),
    .B2(_01786_),
    .ZN(_01983_));
 MUX2_X1 _24955_ (.A(_01725_),
    .B(_01791_),
    .S(_01793_),
    .Z(_01984_));
 BUF_X4 _24956_ (.A(_01787_),
    .Z(_01985_));
 AOI21_X1 _24957_ (.A(_01983_),
    .B1(_01984_),
    .B2(_01985_),
    .ZN(_01986_));
 AOI21_X1 _24958_ (.A(_15106_),
    .B1(_01752_),
    .B2(_01914_),
    .ZN(_01987_));
 OAI21_X1 _24959_ (.A(_01848_),
    .B1(_01722_),
    .B2(net523),
    .ZN(_01988_));
 OAI221_X2 _24960_ (.A(_01965_),
    .B1(_01800_),
    .B2(_01986_),
    .C1(_01987_),
    .C2(_01988_),
    .ZN(_01989_));
 NOR2_X1 _24961_ (.A1(_01799_),
    .A2(_01704_),
    .ZN(_01990_));
 OR2_X1 _24962_ (.A1(_01823_),
    .A2(_01884_),
    .ZN(_01991_));
 OAI221_X1 _24963_ (.A(_01990_),
    .B1(_01991_),
    .B2(net757),
    .C1(_01715_),
    .C2(_01701_),
    .ZN(_01992_));
 AND3_X1 _24964_ (.A1(_01842_),
    .A2(_01850_),
    .A3(_01950_),
    .ZN(_01993_));
 NOR3_X2 _24965_ (.A1(net761),
    .A2(_01754_),
    .A3(_01755_),
    .ZN(_01994_));
 AOI21_X1 _24966_ (.A(_01994_),
    .B1(_01977_),
    .B2(_15092_),
    .ZN(_01995_));
 AOI21_X1 _24967_ (.A(_01993_),
    .B1(_01995_),
    .B2(_15106_),
    .ZN(_01996_));
 OAI21_X1 _24968_ (.A(_01992_),
    .B1(_01996_),
    .B2(_01853_),
    .ZN(_01997_));
 OAI21_X1 _24969_ (.A(_01735_),
    .B1(_01989_),
    .B2(_01997_),
    .ZN(_01998_));
 OAI221_X2 _24970_ (.A(_01948_),
    .B1(_01963_),
    .B2(_01964_),
    .C1(_01982_),
    .C2(_01998_),
    .ZN(_00106_));
 NOR2_X1 _24971_ (.A1(_01807_),
    .A2(_01808_),
    .ZN(_01999_));
 NAND2_X2 _24972_ (.A1(_01652_),
    .A2(_01830_),
    .ZN(_02000_));
 NOR3_X2 _24973_ (.A1(_01789_),
    .A2(_01754_),
    .A3(_01755_),
    .ZN(_02001_));
 NOR3_X1 _24974_ (.A1(_01985_),
    .A2(_01971_),
    .A3(_02001_),
    .ZN(_02002_));
 NAND2_X1 _24975_ (.A1(net1201),
    .A2(_01768_),
    .ZN(_02003_));
 AOI21_X2 _24976_ (.A(_01897_),
    .B1(_01895_),
    .B2(_02003_),
    .ZN(_02004_));
 NOR2_X1 _24977_ (.A1(_01747_),
    .A2(_01783_),
    .ZN(_02005_));
 AND2_X1 _24978_ (.A1(_15097_),
    .A2(_01782_),
    .ZN(_02006_));
 OAI33_X1 _24979_ (.A1(_02000_),
    .A2(_02002_),
    .A3(_02004_),
    .B1(_02005_),
    .B2(_02006_),
    .B3(_01764_),
    .ZN(_02007_));
 NAND2_X1 _24980_ (.A1(_01725_),
    .A2(_01769_),
    .ZN(_02008_));
 NAND3_X1 _24981_ (.A1(_01791_),
    .A2(_01651_),
    .A3(_01700_),
    .ZN(_02009_));
 AOI21_X1 _24982_ (.A(_01985_),
    .B1(_02008_),
    .B2(_02009_),
    .ZN(_02010_));
 NOR3_X1 _24983_ (.A1(net1133),
    .A2(_01797_),
    .A3(_01758_),
    .ZN(_02011_));
 NAND3_X1 _24984_ (.A1(_01838_),
    .A2(_01799_),
    .A3(_01700_),
    .ZN(_02012_));
 NAND3_X1 _24985_ (.A1(_01637_),
    .A2(_01651_),
    .A3(_01823_),
    .ZN(_02013_));
 AOI21_X1 _24986_ (.A(_01789_),
    .B1(_02012_),
    .B2(_02013_),
    .ZN(_02014_));
 NOR4_X1 _24987_ (.A1(_01729_),
    .A2(_02010_),
    .A3(_02011_),
    .A4(_02014_),
    .ZN(_02015_));
 OAI21_X1 _24988_ (.A(_01999_),
    .B1(_02007_),
    .B2(_02015_),
    .ZN(_02016_));
 AOI21_X1 _24989_ (.A(_01663_),
    .B1(_01740_),
    .B2(_01803_),
    .ZN(_02017_));
 AOI221_X2 _24990_ (.A(_01823_),
    .B1(_01704_),
    .B2(_01791_),
    .C1(_15097_),
    .C2(_01838_),
    .ZN(_02018_));
 AOI21_X1 _24991_ (.A(_15106_),
    .B1(_01729_),
    .B2(_15086_),
    .ZN(_02019_));
 OAI21_X1 _24992_ (.A(_02018_),
    .B1(_02019_),
    .B2(net126),
    .ZN(_02020_));
 XNOR2_X1 _24993_ (.A(_01897_),
    .B(_01739_),
    .ZN(_02021_));
 OAI21_X4 _24994_ (.A(_01635_),
    .B1(_01670_),
    .B2(_01674_),
    .ZN(_02022_));
 OAI221_X1 _24995_ (.A(_01801_),
    .B1(_02021_),
    .B2(net806),
    .C1(_02022_),
    .C2(_15092_),
    .ZN(_02023_));
 NAND3_X1 _24996_ (.A1(_02017_),
    .A2(_02020_),
    .A3(_02023_),
    .ZN(_02024_));
 AND3_X1 _24997_ (.A1(_01743_),
    .A2(_01651_),
    .A3(_01957_),
    .ZN(_02025_));
 NOR2_X1 _24998_ (.A1(_01799_),
    .A2(_02001_),
    .ZN(_02026_));
 AOI221_X2 _24999_ (.A(_01728_),
    .B1(_02003_),
    .B2(_02025_),
    .C1(_02026_),
    .C2(_01960_),
    .ZN(_02027_));
 MUX2_X1 _25000_ (.A(_01774_),
    .B(_01941_),
    .S(_01636_),
    .Z(_02028_));
 MUX2_X1 _25001_ (.A(_01804_),
    .B(_02028_),
    .S(_01724_),
    .Z(_02029_));
 OAI21_X4 _25002_ (.A(_02027_),
    .B1(_02029_),
    .B2(_01732_),
    .ZN(_02030_));
 AOI21_X1 _25003_ (.A(_01803_),
    .B1(_15086_),
    .B2(net763),
    .ZN(_02031_));
 OAI221_X1 _25004_ (.A(_01990_),
    .B1(_02031_),
    .B2(_01769_),
    .C1(_01745_),
    .C2(_01714_),
    .ZN(_02032_));
 NOR3_X4 _25005_ (.A1(_01774_),
    .A2(_01754_),
    .A3(_01755_),
    .ZN(_02033_));
 NOR3_X2 _25006_ (.A1(_02033_),
    .A2(_01741_),
    .A3(_01639_),
    .ZN(_02034_));
 NAND3_X1 _25007_ (.A1(_01771_),
    .A2(_01685_),
    .A3(_01690_),
    .ZN(_02035_));
 AOI21_X1 _25008_ (.A(_01636_),
    .B1(_01820_),
    .B2(_02035_),
    .ZN(_02036_));
 OR3_X2 _25009_ (.A1(_02034_),
    .A2(_01764_),
    .A3(_02036_),
    .ZN(_02037_));
 AND3_X4 _25010_ (.A1(_01861_),
    .A2(_02032_),
    .A3(_02037_),
    .ZN(_02038_));
 AOI21_X2 _25011_ (.A(_01718_),
    .B1(_01685_),
    .B2(_01690_),
    .ZN(_02039_));
 NOR3_X1 _25012_ (.A1(_01759_),
    .A2(_01754_),
    .A3(_01755_),
    .ZN(_02040_));
 NOR3_X1 _25013_ (.A1(_01842_),
    .A2(_02039_),
    .A3(_02040_),
    .ZN(_02041_));
 NOR3_X1 _25014_ (.A1(_01897_),
    .A2(_01871_),
    .A3(net1130),
    .ZN(_02042_));
 OAI21_X1 _25015_ (.A(_01705_),
    .B1(_02041_),
    .B2(_02042_),
    .ZN(_02043_));
 NAND3_X1 _25016_ (.A1(_01897_),
    .A2(_01786_),
    .A3(_01845_),
    .ZN(_02044_));
 AOI21_X1 _25017_ (.A(_01872_),
    .B1(_01724_),
    .B2(_15092_),
    .ZN(_02045_));
 OAI21_X1 _25018_ (.A(_02044_),
    .B1(_02045_),
    .B2(_15106_),
    .ZN(_02046_));
 OAI21_X1 _25019_ (.A(_02043_),
    .B1(_02046_),
    .B2(_01740_),
    .ZN(_02047_));
 AOI22_X4 _25020_ (.A1(_02038_),
    .A2(_02030_),
    .B1(_02047_),
    .B2(_01738_),
    .ZN(_02048_));
 INV_X1 _25021_ (.A(_01964_),
    .ZN(_02049_));
 AOI21_X1 _25022_ (.A(_15086_),
    .B1(_01897_),
    .B2(_01794_),
    .ZN(_02050_));
 OAI22_X1 _25023_ (.A1(_01718_),
    .A2(_01722_),
    .B1(_01758_),
    .B2(net126),
    .ZN(_02051_));
 NOR3_X1 _25024_ (.A1(_01652_),
    .A2(_02050_),
    .A3(_02051_),
    .ZN(_02052_));
 NAND2_X1 _25025_ (.A1(_01746_),
    .A2(_01743_),
    .ZN(_02053_));
 NAND2_X1 _25026_ (.A1(_01639_),
    .A2(_01970_),
    .ZN(_02054_));
 AOI21_X2 _25027_ (.A(_01699_),
    .B1(_02053_),
    .B2(_02054_),
    .ZN(_02055_));
 NOR3_X2 _25028_ (.A1(_01797_),
    .A2(_01923_),
    .A3(_02055_),
    .ZN(_02056_));
 OR2_X2 _25029_ (.A1(_01705_),
    .A2(_02056_),
    .ZN(_02057_));
 AOI221_X2 _25030_ (.A(_01750_),
    .B1(_01799_),
    .B2(_01723_),
    .C1(_01793_),
    .C2(_01844_),
    .ZN(_02058_));
 AOI21_X1 _25031_ (.A(_01985_),
    .B1(_01652_),
    .B2(_01892_),
    .ZN(_02059_));
 OAI21_X2 _25032_ (.A(_01746_),
    .B1(_01719_),
    .B2(_01720_),
    .ZN(_02060_));
 AND2_X4 _25033_ (.A1(_01786_),
    .A2(_02060_),
    .ZN(_02061_));
 NAND2_X1 _25034_ (.A1(_01798_),
    .A2(_02061_),
    .ZN(_02062_));
 AOI21_X1 _25035_ (.A(_02058_),
    .B1(_02059_),
    .B2(_02062_),
    .ZN(_02063_));
 OAI221_X2 _25036_ (.A(_02049_),
    .B1(_02057_),
    .B2(_02052_),
    .C1(_02063_),
    .C2(_01729_),
    .ZN(_02064_));
 AND4_X4 _25037_ (.A1(_02048_),
    .A2(_02024_),
    .A3(_02016_),
    .A4(_02064_),
    .ZN(_00107_));
 NAND2_X1 _25038_ (.A1(_01809_),
    .A2(_01704_),
    .ZN(_02065_));
 NAND3_X4 _25039_ (.A1(_01950_),
    .A2(_01850_),
    .A3(_01713_),
    .ZN(_02066_));
 AOI21_X4 _25040_ (.A(_01772_),
    .B1(_02066_),
    .B2(_02065_),
    .ZN(_02067_));
 NOR3_X2 _25041_ (.A1(net761),
    .A2(_01744_),
    .A3(_01713_),
    .ZN(_02068_));
 XNOR2_X1 _25042_ (.A(_01744_),
    .B(_01703_),
    .ZN(_02069_));
 NOR2_X1 _25043_ (.A1(_01792_),
    .A2(_01703_),
    .ZN(_02070_));
 AOI221_X2 _25044_ (.A(_02068_),
    .B1(_02069_),
    .B2(_01774_),
    .C1(_01747_),
    .C2(_02070_),
    .ZN(_02071_));
 AOI211_X2 _25045_ (.A(_02067_),
    .B(_01652_),
    .C1(_02071_),
    .C2(_01985_),
    .ZN(_02072_));
 AOI21_X1 _25046_ (.A(_01787_),
    .B1(_01816_),
    .B2(_01850_),
    .ZN(_02073_));
 OAI21_X1 _25047_ (.A(_01950_),
    .B1(_01792_),
    .B2(net763),
    .ZN(_02074_));
 AOI21_X1 _25048_ (.A(_02073_),
    .B1(_02074_),
    .B2(_01985_),
    .ZN(_02075_));
 NOR2_X1 _25049_ (.A1(_01769_),
    .A2(_01715_),
    .ZN(_02076_));
 AOI21_X2 _25050_ (.A(_01639_),
    .B1(_01880_),
    .B2(_01883_),
    .ZN(_02077_));
 AOI21_X1 _25051_ (.A(_02077_),
    .B1(_01897_),
    .B2(_01784_),
    .ZN(_02078_));
 AOI21_X1 _25052_ (.A(_02076_),
    .B1(_02078_),
    .B2(_01977_),
    .ZN(_02079_));
 OAI221_X1 _25053_ (.A(_01808_),
    .B1(_02075_),
    .B2(_01853_),
    .C1(_02079_),
    .C2(_02000_),
    .ZN(_02080_));
 NAND3_X1 _25054_ (.A1(_01700_),
    .A2(_01765_),
    .A3(_01824_),
    .ZN(_02081_));
 OAI21_X1 _25055_ (.A(_02081_),
    .B1(_01804_),
    .B2(_01724_),
    .ZN(_02082_));
 AOI21_X1 _25056_ (.A(_01901_),
    .B1(net758),
    .B2(_01977_),
    .ZN(_02083_));
 OAI221_X1 _25057_ (.A(_01965_),
    .B1(_02000_),
    .B2(_02082_),
    .C1(_02083_),
    .C2(_01764_),
    .ZN(_02084_));
 MUX2_X1 _25058_ (.A(_01604_),
    .B(_15097_),
    .S(_01768_),
    .Z(_02085_));
 OAI221_X2 _25059_ (.A(_01926_),
    .B1(_02085_),
    .B2(_01637_),
    .C1(_01895_),
    .C2(_15087_),
    .ZN(_02086_));
 AOI21_X1 _25060_ (.A(_01854_),
    .B1(_01823_),
    .B2(_15092_),
    .ZN(_02087_));
 OAI21_X1 _25061_ (.A(_01837_),
    .B1(_02087_),
    .B2(_01985_),
    .ZN(_02088_));
 AOI22_X2 _25062_ (.A1(_01809_),
    .A2(_01781_),
    .B1(_02086_),
    .B2(_02088_),
    .ZN(_02089_));
 OAI22_X1 _25063_ (.A1(_02080_),
    .A2(_02072_),
    .B1(_02084_),
    .B2(_02089_),
    .ZN(_02090_));
 OAI22_X2 _25064_ (.A1(net593),
    .A2(_01602_),
    .B1(_01670_),
    .B2(_01674_),
    .ZN(_02091_));
 OAI221_X1 _25065_ (.A(_01823_),
    .B1(_01728_),
    .B2(_01765_),
    .C1(_02091_),
    .C2(_01637_),
    .ZN(_02092_));
 OR2_X1 _25066_ (.A1(_01823_),
    .A2(_01803_),
    .ZN(_02093_));
 AOI21_X1 _25067_ (.A(_01791_),
    .B1(_15086_),
    .B2(_02022_),
    .ZN(_02094_));
 OAI21_X1 _25068_ (.A(_02092_),
    .B1(_02093_),
    .B2(_02094_),
    .ZN(_02095_));
 NOR2_X1 _25069_ (.A1(_01842_),
    .A2(_01728_),
    .ZN(_02096_));
 OAI21_X1 _25070_ (.A(net126),
    .B1(_01814_),
    .B2(_02096_),
    .ZN(_02097_));
 AOI21_X1 _25071_ (.A(_01965_),
    .B1(_02095_),
    .B2(_02097_),
    .ZN(_02098_));
 OAI22_X1 _25072_ (.A1(_15104_),
    .A2(_01758_),
    .B1(_01892_),
    .B2(_01787_),
    .ZN(_02099_));
 OAI21_X1 _25073_ (.A(_01661_),
    .B1(_01739_),
    .B2(_02099_),
    .ZN(_02100_));
 OAI21_X1 _25074_ (.A(_01838_),
    .B1(_01872_),
    .B2(_01869_),
    .ZN(_02101_));
 OAI21_X1 _25075_ (.A(_02101_),
    .B1(_01927_),
    .B2(_01897_),
    .ZN(_02102_));
 AOI21_X1 _25076_ (.A(_02100_),
    .B1(_02102_),
    .B2(_01705_),
    .ZN(_02103_));
 NAND3_X1 _25077_ (.A1(_01637_),
    .A2(_01786_),
    .A3(_01813_),
    .ZN(_02104_));
 NAND2_X1 _25078_ (.A1(_01816_),
    .A2(_01914_),
    .ZN(_02105_));
 OAI21_X1 _25079_ (.A(_02104_),
    .B1(_02105_),
    .B2(_01842_),
    .ZN(_02106_));
 NOR3_X1 _25080_ (.A1(_02106_),
    .A2(_01705_),
    .A3(_01808_),
    .ZN(_02107_));
 OAI21_X2 _25081_ (.A(_01636_),
    .B1(_01792_),
    .B2(_01603_),
    .ZN(_02108_));
 AOI21_X1 _25082_ (.A(_02108_),
    .B1(_01700_),
    .B2(_01718_),
    .ZN(_02109_));
 NOR2_X1 _25083_ (.A1(_01704_),
    .A2(_01803_),
    .ZN(_02110_));
 NAND2_X1 _25084_ (.A1(_01736_),
    .A2(_02110_),
    .ZN(_02111_));
 NAND3_X1 _25085_ (.A1(_01661_),
    .A2(_01739_),
    .A3(_01915_),
    .ZN(_02112_));
 OAI221_X1 _25086_ (.A(_01798_),
    .B1(_02109_),
    .B2(_02111_),
    .C1(_02112_),
    .C2(_15106_),
    .ZN(_02113_));
 NAND2_X1 _25087_ (.A1(_01736_),
    .A2(_01703_),
    .ZN(_02114_));
 AOI221_X2 _25088_ (.A(_02114_),
    .B1(_01909_),
    .B2(_01639_),
    .C1(_01809_),
    .C2(_01768_),
    .ZN(_02115_));
 OAI33_X1 _25089_ (.A1(_02103_),
    .A2(_02098_),
    .A3(_01798_),
    .B1(_02113_),
    .B2(_02107_),
    .B3(_02115_),
    .ZN(_02116_));
 MUX2_X1 _25090_ (.A(_02090_),
    .B(_02116_),
    .S(_01807_),
    .Z(_00108_));
 NAND3_X1 _25091_ (.A1(_01735_),
    .A2(_01786_),
    .A3(_01840_),
    .ZN(_02117_));
 NAND3_X1 _25092_ (.A1(_01900_),
    .A2(_01807_),
    .A3(_01701_),
    .ZN(_02118_));
 AOI21_X1 _25093_ (.A(_15113_),
    .B1(_02117_),
    .B2(_02118_),
    .ZN(_02119_));
 NAND3_X1 _25094_ (.A1(_15113_),
    .A2(_01820_),
    .A3(_01950_),
    .ZN(_02120_));
 NAND2_X1 _25095_ (.A1(_01965_),
    .A2(_02120_),
    .ZN(_02121_));
 MUX2_X1 _25096_ (.A(_01789_),
    .B(_01725_),
    .S(_01792_),
    .Z(_02122_));
 AOI221_X1 _25097_ (.A(_01656_),
    .B1(_01782_),
    .B2(_01791_),
    .C1(_02122_),
    .C2(_01842_),
    .ZN(_02123_));
 OAI21_X1 _25098_ (.A(_15106_),
    .B1(_01801_),
    .B2(_01815_),
    .ZN(_02124_));
 NAND2_X1 _25099_ (.A1(_01850_),
    .A2(_02124_),
    .ZN(_02125_));
 AOI21_X1 _25100_ (.A(_02123_),
    .B1(_02125_),
    .B2(_01807_),
    .ZN(_02126_));
 OAI221_X2 _25101_ (.A(_01926_),
    .B1(_02119_),
    .B2(_02121_),
    .C1(_02126_),
    .C2(_01965_),
    .ZN(_02127_));
 NAND2_X1 _25102_ (.A1(_01750_),
    .A2(_02061_),
    .ZN(_02128_));
 AOI21_X1 _25103_ (.A(_01734_),
    .B1(_01723_),
    .B2(_01636_),
    .ZN(_02129_));
 OAI21_X1 _25104_ (.A(_01636_),
    .B1(_01912_),
    .B2(_02039_),
    .ZN(_02130_));
 OAI21_X1 _25105_ (.A(_02130_),
    .B1(_01721_),
    .B2(net806),
    .ZN(_02131_));
 AOI221_X1 _25106_ (.A(_01661_),
    .B1(_02128_),
    .B2(_02129_),
    .C1(_02131_),
    .C2(_01734_),
    .ZN(_02132_));
 NAND2_X1 _25107_ (.A1(_01771_),
    .A2(_01782_),
    .ZN(_02133_));
 AND2_X1 _25108_ (.A1(_01734_),
    .A2(_01820_),
    .ZN(_02134_));
 OAI22_X1 _25109_ (.A1(_01900_),
    .A2(_01721_),
    .B1(_01758_),
    .B2(_01826_),
    .ZN(_02135_));
 AOI21_X1 _25110_ (.A(_02135_),
    .B1(_01783_),
    .B2(_15086_),
    .ZN(_02136_));
 AOI221_X1 _25111_ (.A(_01736_),
    .B1(_02133_),
    .B2(_02134_),
    .C1(_02136_),
    .C2(_01656_),
    .ZN(_02137_));
 OR3_X2 _25112_ (.A1(_02000_),
    .A2(_02132_),
    .A3(_02137_),
    .ZN(_02138_));
 NAND2_X1 _25113_ (.A1(_01844_),
    .A2(_01637_),
    .ZN(_02139_));
 AOI221_X2 _25114_ (.A(_01728_),
    .B1(_01969_),
    .B2(net761),
    .C1(_02139_),
    .C2(_01769_),
    .ZN(_02140_));
 OAI21_X2 _25115_ (.A(_15106_),
    .B1(_01971_),
    .B2(_01901_),
    .ZN(_02141_));
 AOI21_X2 _25116_ (.A(_01705_),
    .B1(_02141_),
    .B2(_01979_),
    .ZN(_02142_));
 OAI21_X2 _25117_ (.A(_01965_),
    .B1(_02142_),
    .B2(_02140_),
    .ZN(_02143_));
 NAND2_X1 _25118_ (.A1(_15113_),
    .A2(_01892_),
    .ZN(_02144_));
 NOR3_X2 _25119_ (.A1(_01724_),
    .A2(_01830_),
    .A3(_01922_),
    .ZN(_02145_));
 NOR2_X1 _25120_ (.A1(_01871_),
    .A2(_02091_),
    .ZN(_02146_));
 NOR2_X1 _25121_ (.A1(_02145_),
    .A2(_02146_),
    .ZN(_02147_));
 NOR2_X1 _25122_ (.A1(_15092_),
    .A2(_02022_),
    .ZN(_02148_));
 NOR3_X1 _25123_ (.A1(net126),
    .A2(_15086_),
    .A3(_01728_),
    .ZN(_02149_));
 OAI21_X1 _25124_ (.A(_01701_),
    .B1(_02148_),
    .B2(_02149_),
    .ZN(_02150_));
 NAND4_X1 _25125_ (.A1(_01808_),
    .A2(_02144_),
    .A3(_02147_),
    .A4(_02150_),
    .ZN(_02151_));
 NAND4_X1 _25126_ (.A1(_02143_),
    .A2(_01735_),
    .A3(_01798_),
    .A4(_02151_),
    .ZN(_02152_));
 NOR2_X1 _25127_ (.A1(_01768_),
    .A2(_02053_),
    .ZN(_02153_));
 NOR4_X2 _25128_ (.A1(_01757_),
    .A2(_01872_),
    .A3(_02114_),
    .A4(_02153_),
    .ZN(_02154_));
 NAND2_X1 _25129_ (.A1(_15097_),
    .A2(_01782_),
    .ZN(_02155_));
 OAI21_X1 _25130_ (.A(_01802_),
    .B1(_01768_),
    .B2(net125),
    .ZN(_02156_));
 AOI221_X2 _25131_ (.A(_01736_),
    .B1(_01711_),
    .B2(_01712_),
    .C1(_02155_),
    .C2(_02156_),
    .ZN(_02157_));
 NOR4_X2 _25132_ (.A1(_02154_),
    .A2(_01735_),
    .A3(_01732_),
    .A4(_02157_),
    .ZN(_02158_));
 MUX2_X1 _25133_ (.A(_01844_),
    .B(_01815_),
    .S(_01640_),
    .Z(_02159_));
 OAI221_X2 _25134_ (.A(_01832_),
    .B1(_02159_),
    .B2(_01701_),
    .C1(_01670_),
    .C2(_01674_),
    .ZN(_02160_));
 AOI21_X1 _25135_ (.A(net1131),
    .B1(_01701_),
    .B2(net126),
    .ZN(_02161_));
 OAI21_X1 _25136_ (.A(_01957_),
    .B1(_01701_),
    .B2(_01751_),
    .ZN(_02162_));
 MUX2_X1 _25137_ (.A(_02161_),
    .B(_02162_),
    .S(_15113_),
    .Z(_02163_));
 NAND2_X1 _25138_ (.A1(_01965_),
    .A2(_01740_),
    .ZN(_02164_));
 OAI221_X2 _25139_ (.A(_02158_),
    .B1(_02160_),
    .B2(_01965_),
    .C1(_02163_),
    .C2(_02164_),
    .ZN(_02165_));
 NAND4_X1 _25140_ (.A1(_02127_),
    .A2(_02152_),
    .A3(_02165_),
    .A4(_02138_),
    .ZN(_00109_));
 NOR2_X1 _25141_ (.A1(_01734_),
    .A2(_01830_),
    .ZN(_02166_));
 AOI21_X1 _25142_ (.A(_01869_),
    .B1(_01769_),
    .B2(_01809_),
    .ZN(_02167_));
 OAI221_X1 _25143_ (.A(_02166_),
    .B1(_02167_),
    .B2(_01985_),
    .C1(_01753_),
    .C2(_01745_),
    .ZN(_02168_));
 NAND2_X1 _25144_ (.A1(_01774_),
    .A2(_01699_),
    .ZN(_02169_));
 AOI221_X2 _25145_ (.A(_01704_),
    .B1(_02169_),
    .B2(_01960_),
    .C1(_01742_),
    .C2(_01772_),
    .ZN(_02170_));
 MUX2_X1 _25146_ (.A(_01774_),
    .B(_01751_),
    .S(_01635_),
    .Z(_02171_));
 MUX2_X1 _25147_ (.A(_15109_),
    .B(_02171_),
    .S(_01793_),
    .Z(_02172_));
 OAI21_X2 _25148_ (.A(_01735_),
    .B1(_02172_),
    .B2(_01830_),
    .ZN(_02173_));
 NOR2_X1 _25149_ (.A1(_01734_),
    .A2(_01739_),
    .ZN(_02174_));
 INV_X1 _25150_ (.A(_02174_),
    .ZN(_02175_));
 NOR3_X1 _25151_ (.A1(_15107_),
    .A2(_15116_),
    .A3(_01769_),
    .ZN(_02176_));
 MUX2_X1 _25152_ (.A(_15086_),
    .B(_01772_),
    .S(_01791_),
    .Z(_02177_));
 AOI21_X1 _25153_ (.A(_02176_),
    .B1(_02177_),
    .B2(_01801_),
    .ZN(_02178_));
 OAI221_X2 _25154_ (.A(_02168_),
    .B1(_02173_),
    .B2(_02170_),
    .C1(_02175_),
    .C2(_02178_),
    .ZN(_02179_));
 NAND3_X2 _25155_ (.A1(_02179_),
    .A2(_01808_),
    .A3(_01798_),
    .ZN(_02180_));
 OAI21_X1 _25156_ (.A(_01830_),
    .B1(_01715_),
    .B2(_01724_),
    .ZN(_02181_));
 MUX2_X1 _25157_ (.A(_01751_),
    .B(_01802_),
    .S(_01638_),
    .Z(_02182_));
 MUX2_X1 _25158_ (.A(_15118_),
    .B(_02182_),
    .S(_01793_),
    .Z(_02183_));
 AOI22_X2 _25159_ (.A1(_01735_),
    .A2(_02181_),
    .B1(_02183_),
    .B2(_01705_),
    .ZN(_02184_));
 NOR2_X1 _25160_ (.A1(_01733_),
    .A2(_02022_),
    .ZN(_02185_));
 NOR3_X1 _25161_ (.A1(_01636_),
    .A2(_01734_),
    .A3(_01703_),
    .ZN(_02186_));
 AOI221_X2 _25162_ (.A(_01736_),
    .B1(_01813_),
    .B2(_02185_),
    .C1(_02186_),
    .C2(_02061_),
    .ZN(_02187_));
 NOR2_X1 _25163_ (.A1(_15092_),
    .A2(_01722_),
    .ZN(_02188_));
 NOR3_X1 _25164_ (.A1(_01830_),
    .A2(_01778_),
    .A3(_02188_),
    .ZN(_02189_));
 NOR2_X1 _25165_ (.A1(_01809_),
    .A2(_01724_),
    .ZN(_02190_));
 NOR2_X1 _25166_ (.A1(_01941_),
    .A2(_01823_),
    .ZN(_02191_));
 OAI21_X1 _25167_ (.A(_01985_),
    .B1(_02190_),
    .B2(_02191_),
    .ZN(_02192_));
 AOI22_X2 _25168_ (.A1(_02187_),
    .A2(_02184_),
    .B1(_02189_),
    .B2(_02192_),
    .ZN(_02193_));
 NAND3_X1 _25169_ (.A1(_01977_),
    .A2(_01773_),
    .A3(_01824_),
    .ZN(_02194_));
 MUX2_X1 _25170_ (.A(net1201),
    .B(_01809_),
    .S(_01636_),
    .Z(_02195_));
 NAND2_X1 _25171_ (.A1(_01701_),
    .A2(_02195_),
    .ZN(_02196_));
 NAND3_X1 _25172_ (.A1(_02174_),
    .A2(_02194_),
    .A3(_02196_),
    .ZN(_02197_));
 NOR2_X1 _25173_ (.A1(_01807_),
    .A2(_01830_),
    .ZN(_02198_));
 OAI221_X1 _25174_ (.A(_02198_),
    .B1(_02191_),
    .B2(_02108_),
    .C1(_01751_),
    .C2(_01722_),
    .ZN(_02199_));
 NAND3_X1 _25175_ (.A1(_01808_),
    .A2(_02197_),
    .A3(_02199_),
    .ZN(_02200_));
 NAND2_X1 _25176_ (.A1(_01807_),
    .A2(_01705_),
    .ZN(_02201_));
 AND3_X1 _25177_ (.A1(_01640_),
    .A2(_01839_),
    .A3(_02060_),
    .ZN(_02202_));
 AOI21_X1 _25178_ (.A(_02001_),
    .B1(_01970_),
    .B2(_01977_),
    .ZN(_02203_));
 AOI21_X2 _25179_ (.A(_02202_),
    .B1(_02203_),
    .B2(_15113_),
    .ZN(_02204_));
 AOI21_X1 _25180_ (.A(_01838_),
    .B1(_01865_),
    .B2(_01786_),
    .ZN(_02205_));
 AOI21_X1 _25181_ (.A(_01741_),
    .B1(_01970_),
    .B2(_01724_),
    .ZN(_02206_));
 AOI21_X2 _25182_ (.A(_02205_),
    .B1(_02206_),
    .B2(_15106_),
    .ZN(_02207_));
 NAND2_X1 _25183_ (.A1(_01735_),
    .A2(_01729_),
    .ZN(_02208_));
 OAI22_X2 _25184_ (.A1(_02201_),
    .A2(_02204_),
    .B1(_02207_),
    .B2(_02208_),
    .ZN(_02209_));
 OAI211_X2 _25185_ (.A(_01732_),
    .B(_02193_),
    .C1(_02200_),
    .C2(_02209_),
    .ZN(_02210_));
 NOR4_X2 _25186_ (.A1(net523),
    .A2(_01743_),
    .A3(_01754_),
    .A4(_01755_),
    .ZN(_02211_));
 NOR4_X2 _25187_ (.A1(_01734_),
    .A2(_01728_),
    .A3(_01833_),
    .A4(_02211_),
    .ZN(_02212_));
 AOI21_X1 _25188_ (.A(_02212_),
    .B1(_02185_),
    .B2(_01752_),
    .ZN(_02213_));
 AOI21_X1 _25189_ (.A(_01813_),
    .B1(_02212_),
    .B2(_15092_),
    .ZN(_02214_));
 OR2_X1 _25190_ (.A1(_02213_),
    .A2(_02214_),
    .ZN(_02215_));
 AND2_X1 _25191_ (.A1(_01793_),
    .A2(_02053_),
    .ZN(_02216_));
 AOI22_X2 _25192_ (.A1(_15108_),
    .A2(_01977_),
    .B1(_01966_),
    .B2(_02216_),
    .ZN(_02217_));
 OAI21_X1 _25193_ (.A(_01705_),
    .B1(_01722_),
    .B2(net806),
    .ZN(_02218_));
 OAI221_X1 _25194_ (.A(_01735_),
    .B1(_01740_),
    .B2(_02217_),
    .C1(_02218_),
    .C2(_02004_),
    .ZN(_02219_));
 NAND2_X1 _25195_ (.A1(_01801_),
    .A2(_01803_),
    .ZN(_02220_));
 NAND4_X1 _25196_ (.A1(net126),
    .A2(_01979_),
    .A3(_02174_),
    .A4(_02220_),
    .ZN(_02221_));
 NOR2_X1 _25197_ (.A1(_01732_),
    .A2(_01808_),
    .ZN(_02222_));
 NAND4_X1 _25198_ (.A1(_02215_),
    .A2(_02219_),
    .A3(_02221_),
    .A4(_02222_),
    .ZN(_02223_));
 AND3_X4 _25199_ (.A1(_02180_),
    .A2(_02210_),
    .A3(_02223_),
    .ZN(_00110_));
 NAND3_X1 _25200_ (.A1(_01732_),
    .A2(_01807_),
    .A3(_01965_),
    .ZN(_02224_));
 OAI221_X1 _25201_ (.A(_02144_),
    .B1(_01722_),
    .B2(net1201),
    .C1(net806),
    .C2(_01973_),
    .ZN(_02225_));
 OAI21_X1 _25202_ (.A(_01740_),
    .B1(_02224_),
    .B2(_02225_),
    .ZN(_02226_));
 OAI221_X1 _25203_ (.A(_01798_),
    .B1(_01701_),
    .B2(_01771_),
    .C1(_01758_),
    .C2(_01753_),
    .ZN(_02227_));
 NAND2_X1 _25204_ (.A1(_01662_),
    .A2(_02227_),
    .ZN(_02228_));
 NOR2_X1 _25205_ (.A1(_01809_),
    .A2(_01842_),
    .ZN(_02229_));
 NOR3_X1 _25206_ (.A1(_01801_),
    .A2(net757),
    .A3(_02229_),
    .ZN(_02230_));
 AOI21_X1 _25207_ (.A(_02230_),
    .B1(_01801_),
    .B2(_15116_),
    .ZN(_02231_));
 AOI21_X1 _25208_ (.A(_02228_),
    .B1(_02231_),
    .B2(_01732_),
    .ZN(_02232_));
 AOI21_X1 _25209_ (.A(_01740_),
    .B1(_02195_),
    .B2(_01701_),
    .ZN(_02233_));
 OAI21_X1 _25210_ (.A(_01801_),
    .B1(_01803_),
    .B2(_02077_),
    .ZN(_02234_));
 AOI21_X1 _25211_ (.A(_02224_),
    .B1(_02233_),
    .B2(_02234_),
    .ZN(_02235_));
 OAI21_X1 _25212_ (.A(_02226_),
    .B1(_02232_),
    .B2(_02235_),
    .ZN(_02236_));
 NOR2_X1 _25213_ (.A1(_01725_),
    .A2(_01977_),
    .ZN(_02237_));
 OAI221_X1 _25214_ (.A(_01990_),
    .B1(_02108_),
    .B2(_02237_),
    .C1(_15113_),
    .C2(_01718_),
    .ZN(_02238_));
 AND2_X1 _25215_ (.A1(_01861_),
    .A2(_02238_),
    .ZN(_02239_));
 AOI21_X1 _25216_ (.A(_01994_),
    .B1(_02177_),
    .B2(_01801_),
    .ZN(_02240_));
 NAND3_X1 _25217_ (.A1(_01985_),
    .A2(_01820_),
    .A3(_02035_),
    .ZN(_02241_));
 AND3_X1 _25218_ (.A1(_01729_),
    .A2(_01870_),
    .A3(_02241_),
    .ZN(_02242_));
 AOI211_X2 _25219_ (.A(_01787_),
    .B(_01971_),
    .C1(_01700_),
    .C2(net763),
    .ZN(_02243_));
 OAI21_X1 _25220_ (.A(_02060_),
    .B1(_01977_),
    .B2(_01771_),
    .ZN(_02244_));
 AOI21_X1 _25221_ (.A(_02243_),
    .B1(_02244_),
    .B2(_15113_),
    .ZN(_02245_));
 AOI21_X1 _25222_ (.A(_02242_),
    .B1(_02245_),
    .B2(_01740_),
    .ZN(_02246_));
 OAI221_X2 _25223_ (.A(_02239_),
    .B1(_02240_),
    .B2(_01853_),
    .C1(_02246_),
    .C2(_01732_),
    .ZN(_02247_));
 NOR2_X1 _25224_ (.A1(_01771_),
    .A2(_01703_),
    .ZN(_02248_));
 NOR2_X1 _25225_ (.A1(_15097_),
    .A2(_01787_),
    .ZN(_02249_));
 AOI221_X2 _25226_ (.A(_01651_),
    .B1(_01969_),
    .B2(_02248_),
    .C1(_02249_),
    .C2(_01691_),
    .ZN(_02250_));
 NOR2_X1 _25227_ (.A1(_01977_),
    .A2(_01728_),
    .ZN(_02251_));
 AOI21_X1 _25228_ (.A(_02251_),
    .B1(_02070_),
    .B2(net126),
    .ZN(_02252_));
 AOI21_X1 _25229_ (.A(_01781_),
    .B1(_01782_),
    .B2(_01729_),
    .ZN(_02253_));
 OAI221_X2 _25230_ (.A(_02250_),
    .B1(_02252_),
    .B2(_15086_),
    .C1(_02253_),
    .C2(net126),
    .ZN(_02254_));
 AOI21_X1 _25231_ (.A(_01969_),
    .B1(_01728_),
    .B2(_01769_),
    .ZN(_02255_));
 AOI21_X1 _25232_ (.A(_02033_),
    .B1(_01691_),
    .B2(_01751_),
    .ZN(_02256_));
 OAI221_X1 _25233_ (.A(_02022_),
    .B1(_02255_),
    .B2(_01900_),
    .C1(_02256_),
    .C2(_15113_),
    .ZN(_02257_));
 AOI21_X1 _25234_ (.A(_01778_),
    .B1(_02257_),
    .B2(_01732_),
    .ZN(_02258_));
 AOI221_X1 _25235_ (.A(_01703_),
    .B1(_01781_),
    .B2(_01747_),
    .C1(_02074_),
    .C2(_01750_),
    .ZN(_02259_));
 AOI21_X1 _25236_ (.A(_01640_),
    .B1(_01839_),
    .B2(_01914_),
    .ZN(_02260_));
 NOR3_X1 _25237_ (.A1(_01637_),
    .A2(_01854_),
    .A3(_02039_),
    .ZN(_02261_));
 NOR3_X1 _25238_ (.A1(_01830_),
    .A2(_02260_),
    .A3(_02261_),
    .ZN(_02262_));
 OR2_X1 _25239_ (.A1(_02259_),
    .A2(_02262_),
    .ZN(_02263_));
 NOR2_X1 _25240_ (.A1(_01732_),
    .A2(_01964_),
    .ZN(_02264_));
 MUX2_X1 _25241_ (.A(_01789_),
    .B(_01603_),
    .S(_01792_),
    .Z(_02265_));
 OAI21_X1 _25242_ (.A(_01908_),
    .B1(_02265_),
    .B2(_01842_),
    .ZN(_02266_));
 OAI21_X2 _25243_ (.A(_01750_),
    .B1(_01872_),
    .B2(_01854_),
    .ZN(_02267_));
 OAI21_X1 _25244_ (.A(_02267_),
    .B1(_01927_),
    .B2(_01897_),
    .ZN(_02268_));
 MUX2_X1 _25245_ (.A(_02266_),
    .B(_02268_),
    .S(_01797_),
    .Z(_02269_));
 NOR2_X1 _25246_ (.A1(_01737_),
    .A2(_01729_),
    .ZN(_02270_));
 AOI222_X2 _25247_ (.A1(_02254_),
    .A2(_02258_),
    .B1(_02263_),
    .B2(_02264_),
    .C1(_02270_),
    .C2(_02269_),
    .ZN(_02271_));
 NAND3_X1 _25248_ (.A1(_02236_),
    .A2(_02247_),
    .A3(_02271_),
    .ZN(_00111_));
 XNOR2_X2 _25249_ (.A(_10503_),
    .B(_10506_),
    .ZN(_02272_));
 XNOR2_X2 _25250_ (.A(_13167_),
    .B(_02272_),
    .ZN(_02273_));
 XOR2_X2 _25251_ (.A(_10453_),
    .B(\sa20_sub[0] ),
    .Z(_02274_));
 XNOR2_X2 _25252_ (.A(_02274_),
    .B(\sa12_sr[1] ),
    .ZN(_02275_));
 XNOR2_X1 _25253_ (.A(_02273_),
    .B(_02275_),
    .ZN(_02276_));
 MUX2_X1 _25254_ (.A(_00470_),
    .B(_02276_),
    .S(_09100_),
    .Z(_02277_));
 XOR2_X2 _25255_ (.A(_06470_),
    .B(_02277_),
    .Z(_02278_));
 INV_X32 _25256_ (.A(net1041),
    .ZN(_02279_));
 BUF_X1 rebuffer219 (.A(_02341_),
    .Z(net724));
 BUF_X4 clone247 (.A(net802),
    .Z(net801));
 XNOR2_X1 _25259_ (.A(net1069),
    .B(net662),
    .ZN(_02281_));
 NAND3_X1 _25260_ (.A1(_06456_),
    .A2(_09099_),
    .A3(_13186_),
    .ZN(_02282_));
 NOR2_X1 _25261_ (.A1(_06456_),
    .A2(_08972_),
    .ZN(_02283_));
 NAND2_X1 _25262_ (.A1(_13179_),
    .A2(_02283_),
    .ZN(_02284_));
 AOI21_X1 _25263_ (.A(_02281_),
    .B1(_02282_),
    .B2(_02284_),
    .ZN(_02285_));
 XOR2_X1 _25264_ (.A(net530),
    .B(_02272_),
    .Z(_02286_));
 NAND2_X1 _25265_ (.A1(_13186_),
    .A2(_02283_),
    .ZN(_02287_));
 NAND3_X1 _25266_ (.A1(_06456_),
    .A2(_09011_),
    .A3(_13179_),
    .ZN(_02288_));
 AOI21_X1 _25267_ (.A(_02286_),
    .B1(_02287_),
    .B2(_02288_),
    .ZN(_02289_));
 INV_X1 _25268_ (.A(_06456_),
    .ZN(_02290_));
 NAND3_X1 _25269_ (.A1(_02290_),
    .A2(_09027_),
    .A3(_00471_),
    .ZN(_02291_));
 NAND2_X1 _25270_ (.A1(_06456_),
    .A2(_09015_),
    .ZN(_02292_));
 OAI21_X1 _25271_ (.A(_02291_),
    .B1(_02292_),
    .B2(_00471_),
    .ZN(_02293_));
 OR3_X2 _25272_ (.A1(_02285_),
    .A2(_02289_),
    .A3(_02293_),
    .ZN(_02294_));
 BUF_X4 _25273_ (.A(_02294_),
    .Z(_02295_));
 INV_X4 _25274_ (.A(_02295_),
    .ZN(_02296_));
 BUF_X8 _25275_ (.A(_02296_),
    .Z(_15133_));
 XOR2_X2 _25276_ (.A(net556),
    .B(_10478_),
    .Z(_02297_));
 XOR2_X2 _25277_ (.A(net545),
    .B(_02297_),
    .Z(_02298_));
 NAND3_X1 _25278_ (.A1(_06482_),
    .A2(_09194_),
    .A3(_13205_),
    .ZN(_02299_));
 NOR2_X1 _25279_ (.A1(_06482_),
    .A2(_09027_),
    .ZN(_02300_));
 NAND2_X1 _25280_ (.A1(_13198_),
    .A2(_02300_),
    .ZN(_02301_));
 AOI21_X2 _25281_ (.A(_02298_),
    .B1(_02299_),
    .B2(_02301_),
    .ZN(_02302_));
 XNOR2_X1 _25282_ (.A(net545),
    .B(_02297_),
    .ZN(_02303_));
 NAND2_X1 _25283_ (.A1(_13205_),
    .A2(_02300_),
    .ZN(_02304_));
 NAND3_X1 _25284_ (.A1(_06482_),
    .A2(_09074_),
    .A3(_13198_),
    .ZN(_02305_));
 AOI21_X2 _25285_ (.A(_02303_),
    .B1(_02304_),
    .B2(_02305_),
    .ZN(_02306_));
 NAND3_X1 _25286_ (.A1(_06489_),
    .A2(_08973_),
    .A3(_00472_),
    .ZN(_02307_));
 NAND2_X1 _25287_ (.A1(_06482_),
    .A2(_08973_),
    .ZN(_02308_));
 OAI21_X2 _25288_ (.A(_02307_),
    .B1(_02308_),
    .B2(_00472_),
    .ZN(_02309_));
 NOR3_X4 _25289_ (.A1(_02302_),
    .A2(_02306_),
    .A3(_02309_),
    .ZN(_02310_));
 INV_X4 _25290_ (.A(net1095),
    .ZN(_02311_));
 BUF_X4 _25291_ (.A(_02311_),
    .Z(_02312_));
 BUF_X4 _25292_ (.A(_02312_),
    .Z(_02313_));
 BUF_X4 _25293_ (.A(_02313_),
    .Z(_15149_));
 BUF_X8 _25294_ (.A(_02278_),
    .Z(_02314_));
 BUF_X2 rebuffer116 (.A(_14862_),
    .Z(net599));
 BUF_X8 _25296_ (.A(_02310_),
    .Z(_02315_));
 BUF_X8 _25297_ (.A(_02315_),
    .Z(_02316_));
 BUF_X4 _25298_ (.A(_02316_),
    .Z(_02317_));
 BUF_X4 _25299_ (.A(_02317_),
    .Z(_02318_));
 BUF_X4 _25300_ (.A(_02318_),
    .Z(_02319_));
 BUF_X8 _25301_ (.A(_02319_),
    .Z(_15142_));
 XNOR2_X1 _25302_ (.A(_10541_),
    .B(_10517_),
    .ZN(_02320_));
 XNOR2_X1 _25303_ (.A(_10536_),
    .B(_10524_),
    .ZN(_02321_));
 XNOR2_X1 _25304_ (.A(_02320_),
    .B(_02321_),
    .ZN(_02322_));
 MUX2_X2 _25305_ (.A(\text_in_r[45] ),
    .B(_02322_),
    .S(_09023_),
    .Z(_02323_));
 XOR2_X2 _25306_ (.A(_06545_),
    .B(_02323_),
    .Z(_02324_));
 BUF_X4 _25307_ (.A(_02324_),
    .Z(_02325_));
 XNOR2_X1 _25308_ (.A(_10512_),
    .B(_10506_),
    .ZN(_02326_));
 XNOR2_X2 _25309_ (.A(_10458_),
    .B(_02326_),
    .ZN(_02327_));
 XNOR2_X1 _25310_ (.A(_10513_),
    .B(_02327_),
    .ZN(_02328_));
 MUX2_X2 _25311_ (.A(\text_in_r[47] ),
    .B(_02328_),
    .S(_09158_),
    .Z(_02329_));
 XOR2_X2 _25312_ (.A(_06567_),
    .B(_02329_),
    .Z(_02330_));
 NAND2_X1 _25313_ (.A1(_02325_),
    .A2(_02330_),
    .ZN(_02331_));
 INV_X2 _25314_ (.A(_15126_),
    .ZN(_02332_));
 BUF_X2 _25315_ (.A(\text_in_r[43] ),
    .Z(_02333_));
 XNOR2_X1 _25316_ (.A(_10535_),
    .B(net712),
    .ZN(_02334_));
 XNOR2_X1 _25317_ (.A(_10475_),
    .B(_10539_),
    .ZN(_02335_));
 XNOR2_X2 _25318_ (.A(_02334_),
    .B(_02335_),
    .ZN(_02336_));
 XNOR2_X1 _25319_ (.A(_10554_),
    .B(_10503_),
    .ZN(_02337_));
 XNOR2_X1 _25320_ (.A(_10479_),
    .B(_02337_),
    .ZN(_02338_));
 XNOR2_X2 _25321_ (.A(_02336_),
    .B(_02338_),
    .ZN(_02339_));
 MUX2_X2 _25322_ (.A(_02333_),
    .B(_02339_),
    .S(_09099_),
    .Z(_02340_));
 XNOR2_X2 _25323_ (.A(_02340_),
    .B(_06516_),
    .ZN(_02341_));
 BUF_X4 _25324_ (.A(net728),
    .Z(_02342_));
 BUF_X4 _25325_ (.A(_02342_),
    .Z(_02343_));
 BUF_X4 _25326_ (.A(_02343_),
    .Z(_02344_));
 NAND2_X1 _25327_ (.A1(_02332_),
    .A2(_02344_),
    .ZN(_02345_));
 BUF_X8 _25328_ (.A(_15129_),
    .Z(_02346_));
 INV_X1 _25329_ (.A(_06516_),
    .ZN(_02347_));
 XNOR2_X2 _25330_ (.A(_02340_),
    .B(_02347_),
    .ZN(_02348_));
 BUF_X4 _25331_ (.A(_02348_),
    .Z(_02349_));
 BUF_X8 _25332_ (.A(_02349_),
    .Z(_02350_));
 NAND2_X1 _25333_ (.A1(_02346_),
    .A2(_02350_),
    .ZN(_02351_));
 NAND3_X1 _25334_ (.A1(_15142_),
    .A2(_02345_),
    .A3(_02351_),
    .ZN(_02352_));
 XNOR2_X1 _25335_ (.A(_10525_),
    .B(_13229_),
    .ZN(_02353_));
 XNOR2_X1 _25336_ (.A(_10502_),
    .B(_02353_),
    .ZN(_02354_));
 MUX2_X2 _25337_ (.A(\text_in_r[46] ),
    .B(_02354_),
    .S(_11191_),
    .Z(_02355_));
 XNOR2_X2 _25338_ (.A(_06558_),
    .B(_02355_),
    .ZN(_02356_));
 XOR2_X2 _25339_ (.A(_10554_),
    .B(net712),
    .Z(_02357_));
 XNOR2_X2 _25340_ (.A(_10528_),
    .B(_02357_),
    .ZN(_02358_));
 XOR2_X1 _25341_ (.A(_13268_),
    .B(_02358_),
    .Z(_02359_));
 MUX2_X2 _25342_ (.A(\text_in_r[44] ),
    .B(_02359_),
    .S(_09075_),
    .Z(_02360_));
 XNOR2_X2 _25343_ (.A(_06532_),
    .B(_02360_),
    .ZN(_02361_));
 BUF_X4 _25344_ (.A(_02361_),
    .Z(_02362_));
 NAND2_X2 _25345_ (.A1(_02356_),
    .A2(_02362_),
    .ZN(_02363_));
 NOR2_X4 _25346_ (.A1(_02315_),
    .A2(net728),
    .ZN(_02364_));
 BUF_X4 split203 (.A(net498),
    .Z(net203));
 CLKBUF_X3 _25348_ (.A(_15136_),
    .Z(_02366_));
 AOI21_X1 _25349_ (.A(_02363_),
    .B1(_02364_),
    .B2(_02366_),
    .ZN(_02367_));
 AOI21_X1 _25350_ (.A(_02331_),
    .B1(_02352_),
    .B2(_02367_),
    .ZN(_02368_));
 XOR2_X2 _25351_ (.A(_06532_),
    .B(_02360_),
    .Z(_02369_));
 NAND2_X2 _25352_ (.A1(_02356_),
    .A2(_02369_),
    .ZN(_02370_));
 CLKBUF_X3 _25353_ (.A(_15134_),
    .Z(_02371_));
 NOR3_X2 _25354_ (.A1(_02371_),
    .A2(_02315_),
    .A3(_02348_),
    .ZN(_02372_));
 OR2_X1 _25355_ (.A1(_02370_),
    .A2(_02372_),
    .ZN(_02373_));
 INV_X2 _25356_ (.A(_15129_),
    .ZN(_02374_));
 BUF_X4 _25357_ (.A(_02342_),
    .Z(_02375_));
 BUF_X4 _25358_ (.A(_02375_),
    .Z(_02376_));
 NAND2_X1 _25359_ (.A1(_02374_),
    .A2(_02376_),
    .ZN(_02377_));
 BUF_X4 _25360_ (.A(_15126_),
    .Z(_02378_));
 BUF_X4 _25361_ (.A(_02349_),
    .Z(_02379_));
 CLKBUF_X3 _25362_ (.A(_02379_),
    .Z(_02380_));
 NAND2_X1 _25363_ (.A1(_02378_),
    .A2(_02380_),
    .ZN(_02381_));
 AOI21_X2 _25364_ (.A(_02313_),
    .B1(_02377_),
    .B2(_02381_),
    .ZN(_02382_));
 BUF_X4 _25365_ (.A(_02369_),
    .Z(_02383_));
 CLKBUF_X3 _25366_ (.A(_02383_),
    .Z(_02384_));
 NOR2_X2 _25367_ (.A1(net731),
    .A2(_02350_),
    .ZN(_02385_));
 NOR2_X4 _25368_ (.A1(_02295_),
    .A2(_02342_),
    .ZN(_02386_));
 NOR3_X1 _25369_ (.A1(_15149_),
    .A2(_02385_),
    .A3(_02386_),
    .ZN(_02387_));
 NOR2_X1 _25370_ (.A1(_02371_),
    .A2(_02344_),
    .ZN(_02388_));
 BUF_X4 _25371_ (.A(_15125_),
    .Z(_02389_));
 BUF_X4 _25372_ (.A(net588),
    .Z(_02390_));
 BUF_X4 _25373_ (.A(_02350_),
    .Z(_02391_));
 NOR2_X2 _25374_ (.A1(_02390_),
    .A2(_02391_),
    .ZN(_02392_));
 NOR3_X1 _25375_ (.A1(_15142_),
    .A2(_02388_),
    .A3(_02392_),
    .ZN(_02393_));
 NOR3_X1 _25376_ (.A1(_02384_),
    .A2(_02387_),
    .A3(_02393_),
    .ZN(_02394_));
 XOR2_X2 _25377_ (.A(_06558_),
    .B(_02355_),
    .Z(_02395_));
 BUF_X4 _25378_ (.A(_02395_),
    .Z(_02396_));
 BUF_X4 _25379_ (.A(_02396_),
    .Z(_02397_));
 TAPCELL_X1 PHY_EDGE_ROW_0_Right_0 ();
 CLKBUF_X3 _25381_ (.A(_15131_),
    .Z(_02399_));
 CLKBUF_X3 _25382_ (.A(_02391_),
    .Z(_02400_));
 MUX2_X1 _25383_ (.A(_02378_),
    .B(_02399_),
    .S(_02400_),
    .Z(_02401_));
 BUF_X4 _25384_ (.A(_02311_),
    .Z(_02402_));
 BUF_X4 _25385_ (.A(net728),
    .Z(_02403_));
 NAND2_X4 _25386_ (.A1(_02402_),
    .A2(_02403_),
    .ZN(_02404_));
 BUF_X4 _25387_ (.A(_15124_),
    .Z(_02405_));
 INV_X1 _25388_ (.A(_02405_),
    .ZN(_02406_));
 BUF_X4 _25389_ (.A(_02406_),
    .Z(_02407_));
 OAI221_X1 _25390_ (.A(_02384_),
    .B1(_02401_),
    .B2(_15149_),
    .C1(_02404_),
    .C2(_02407_),
    .ZN(_02408_));
 NAND2_X1 _25391_ (.A1(_02397_),
    .A2(_02408_),
    .ZN(_02409_));
 OAI221_X2 _25392_ (.A(_02368_),
    .B1(_02373_),
    .B2(_02382_),
    .C1(_02394_),
    .C2(_02409_),
    .ZN(_02410_));
 BUF_X4 _25393_ (.A(_02343_),
    .Z(_02411_));
 MUX2_X1 _25394_ (.A(_02390_),
    .B(_02366_),
    .S(_02411_),
    .Z(_02412_));
 OAI221_X1 _25395_ (.A(_02397_),
    .B1(_02404_),
    .B2(_02399_),
    .C1(_02412_),
    .C2(_15149_),
    .ZN(_02413_));
 BUF_X4 _25396_ (.A(_02356_),
    .Z(_02414_));
 BUF_X4 _25397_ (.A(_02379_),
    .Z(_02415_));
 BUF_X4 _25398_ (.A(_02415_),
    .Z(_02416_));
 AND2_X1 _25399_ (.A1(_15147_),
    .A2(_02416_),
    .ZN(_02417_));
 NAND2_X1 _25400_ (.A1(net588),
    .A2(_02311_),
    .ZN(_02418_));
 NOR2_X1 _25401_ (.A1(_02350_),
    .A2(_02418_),
    .ZN(_02419_));
 OAI21_X1 _25402_ (.A(_02414_),
    .B1(_02417_),
    .B2(_02419_),
    .ZN(_02420_));
 NAND3_X1 _25403_ (.A1(_02384_),
    .A2(_02413_),
    .A3(_02420_),
    .ZN(_02421_));
 INV_X4 _25404_ (.A(net1211),
    .ZN(_02422_));
 MUX2_X1 _25405_ (.A(_02422_),
    .B(_02346_),
    .S(_02315_),
    .Z(_02423_));
 OR2_X4 _25406_ (.A1(_02415_),
    .A2(_02423_),
    .ZN(_02424_));
 NOR2_X2 _25407_ (.A1(_02295_),
    .A2(_02315_),
    .ZN(_02425_));
 CLKBUF_X3 _25408_ (.A(_02312_),
    .Z(_02426_));
 CLKBUF_X3 _25409_ (.A(_02426_),
    .Z(_02427_));
 NOR2_X1 _25410_ (.A1(_02405_),
    .A2(_02427_),
    .ZN(_02428_));
 OAI21_X1 _25411_ (.A(_02416_),
    .B1(_02425_),
    .B2(_02428_),
    .ZN(_02429_));
 NOR2_X2 _25412_ (.A1(_02317_),
    .A2(_02379_),
    .ZN(_02430_));
 AOI21_X1 _25413_ (.A(_02363_),
    .B1(_02430_),
    .B2(_02378_),
    .ZN(_02431_));
 NAND3_X1 _25414_ (.A1(_02424_),
    .A2(_02429_),
    .A3(_02431_),
    .ZN(_02432_));
 XNOR2_X2 _25415_ (.A(_06545_),
    .B(_02323_),
    .ZN(_02433_));
 BUF_X4 _25416_ (.A(_02433_),
    .Z(_02434_));
 BUF_X4 _25417_ (.A(_02434_),
    .Z(_02435_));
 BUF_X4 _25418_ (.A(_02330_),
    .Z(_02436_));
 NAND2_X1 _25419_ (.A1(_02435_),
    .A2(_02436_),
    .ZN(_02437_));
 INV_X1 _25420_ (.A(_02437_),
    .ZN(_02438_));
 NOR2_X2 _25421_ (.A1(_02356_),
    .A2(_02383_),
    .ZN(_02439_));
 BUF_X4 _25422_ (.A(_02344_),
    .Z(_02440_));
 AOI21_X1 _25423_ (.A(_02386_),
    .B1(_02440_),
    .B2(_02399_),
    .ZN(_02441_));
 BUF_X2 _25424_ (.A(_15138_),
    .Z(_02442_));
 CLKBUF_X3 _25425_ (.A(_02442_),
    .Z(_02443_));
 NAND2_X4 _25426_ (.A1(_02315_),
    .A2(net1174),
    .ZN(_02444_));
 OAI221_X2 _25427_ (.A(_02439_),
    .B1(_02441_),
    .B2(_15142_),
    .C1(_02443_),
    .C2(_02444_),
    .ZN(_02445_));
 NAND4_X2 _25428_ (.A1(_02421_),
    .A2(_02432_),
    .A3(_02438_),
    .A4(_02445_),
    .ZN(_02446_));
 BUF_X4 _25429_ (.A(_02325_),
    .Z(_02447_));
 NOR2_X2 _25430_ (.A1(_02447_),
    .A2(_02436_),
    .ZN(_02448_));
 NOR2_X2 _25431_ (.A1(_02356_),
    .A2(_02362_),
    .ZN(_02449_));
 NOR2_X1 _25432_ (.A1(net732),
    .A2(_02416_),
    .ZN(_02450_));
 NOR3_X1 _25433_ (.A1(_15142_),
    .A2(_02386_),
    .A3(_02450_),
    .ZN(_02451_));
 BUF_X4 clone3 (.A(net4),
    .Z(net3));
 INV_X16 _25435_ (.A(net1042),
    .ZN(_02453_));
 NOR2_X2 _25436_ (.A1(_02453_),
    .A2(_02343_),
    .ZN(_02454_));
 NOR2_X2 _25437_ (.A1(net720),
    .A2(_02391_),
    .ZN(_02455_));
 NOR3_X1 _25438_ (.A1(_15149_),
    .A2(_02454_),
    .A3(_02455_),
    .ZN(_02456_));
 OAI21_X1 _25439_ (.A(_02449_),
    .B1(_02451_),
    .B2(_02456_),
    .ZN(_02457_));
 NAND2_X2 _25440_ (.A1(net720),
    .A2(_02312_),
    .ZN(_02458_));
 NOR2_X1 _25441_ (.A1(_06516_),
    .A2(_00991_),
    .ZN(_02459_));
 NAND2_X1 _25442_ (.A1(net506),
    .A2(_02459_),
    .ZN(_02460_));
 NOR2_X1 _25443_ (.A1(_02347_),
    .A2(_00991_),
    .ZN(_02461_));
 NAND2_X1 _25444_ (.A1(_02389_),
    .A2(_02461_),
    .ZN(_02462_));
 MUX2_X1 _25445_ (.A(_02460_),
    .B(_02462_),
    .S(_02339_),
    .Z(_02463_));
 INV_X1 _25446_ (.A(_02333_),
    .ZN(_02464_));
 NAND2_X1 _25447_ (.A1(_02464_),
    .A2(_02389_),
    .ZN(_02465_));
 NAND2_X1 _25448_ (.A1(_02347_),
    .A2(_09823_),
    .ZN(_02466_));
 NAND2_X1 _25449_ (.A1(_06516_),
    .A2(_09823_),
    .ZN(_02467_));
 NAND2_X1 _25450_ (.A1(_02333_),
    .A2(net506),
    .ZN(_02468_));
 OAI22_X2 _25451_ (.A1(_02465_),
    .A2(_02466_),
    .B1(_02467_),
    .B2(_02468_),
    .ZN(_02469_));
 INV_X2 _25452_ (.A(_02469_),
    .ZN(_02470_));
 NAND2_X4 _25453_ (.A1(net1039),
    .A2(_02470_),
    .ZN(_02471_));
 NOR2_X1 _25454_ (.A1(_02390_),
    .A2(_02317_),
    .ZN(_02472_));
 NAND2_X2 _25455_ (.A1(net144),
    .A2(_02375_),
    .ZN(_02473_));
 AOI221_X2 _25456_ (.A(_02370_),
    .B1(_02471_),
    .B2(_02458_),
    .C1(_02472_),
    .C2(_02473_),
    .ZN(_02474_));
 CLKBUF_X3 _25457_ (.A(_02383_),
    .Z(_02475_));
 NAND2_X1 _25458_ (.A1(net1040),
    .A2(_02402_),
    .ZN(_02476_));
 NOR2_X2 _25459_ (.A1(_02378_),
    .A2(_02402_),
    .ZN(_02477_));
 NOR2_X1 _25460_ (.A1(_02415_),
    .A2(_02477_),
    .ZN(_02478_));
 AOI21_X1 _25461_ (.A(_02475_),
    .B1(_02476_),
    .B2(_02478_),
    .ZN(_02479_));
 NOR2_X1 _25462_ (.A1(_02443_),
    .A2(_02312_),
    .ZN(_02480_));
 OAI21_X1 _25463_ (.A(_02380_),
    .B1(_02425_),
    .B2(_02480_),
    .ZN(_02481_));
 AND2_X1 _25464_ (.A1(_02395_),
    .A2(_02481_),
    .ZN(_02482_));
 NOR2_X4 _25465_ (.A1(_02311_),
    .A2(_02341_),
    .ZN(_02483_));
 XNOR2_X2 _25466_ (.A(_02315_),
    .B(net728),
    .ZN(_02484_));
 AOI221_X2 _25467_ (.A(_02372_),
    .B1(_02483_),
    .B2(_02390_),
    .C1(_02484_),
    .C2(_02407_),
    .ZN(_02485_));
 NOR2_X2 _25468_ (.A1(_02396_),
    .A2(_02384_),
    .ZN(_02486_));
 AOI221_X2 _25469_ (.A(_02474_),
    .B1(_02479_),
    .B2(_02482_),
    .C1(_02485_),
    .C2(_02486_),
    .ZN(_02487_));
 NAND3_X2 _25470_ (.A1(_02448_),
    .A2(_02457_),
    .A3(_02487_),
    .ZN(_02488_));
 NOR2_X1 _25471_ (.A1(_02399_),
    .A2(_02444_),
    .ZN(_02489_));
 BUF_X4 _25472_ (.A(_02295_),
    .Z(_15122_));
 NAND2_X1 _25473_ (.A1(_15122_),
    .A2(_02344_),
    .ZN(_02490_));
 AOI21_X1 _25474_ (.A(_15142_),
    .B1(_02351_),
    .B2(_02490_),
    .ZN(_02491_));
 OAI21_X1 _25475_ (.A(_02439_),
    .B1(_02489_),
    .B2(_02491_),
    .ZN(_02492_));
 NOR3_X1 _25476_ (.A1(_15149_),
    .A2(_02388_),
    .A3(_02471_),
    .ZN(_02493_));
 NAND2_X1 _25477_ (.A1(_02407_),
    .A2(_02416_),
    .ZN(_02494_));
 INV_X2 _25478_ (.A(_02442_),
    .ZN(_02495_));
 NAND2_X1 _25479_ (.A1(_02495_),
    .A2(_02411_),
    .ZN(_02496_));
 AND3_X1 _25480_ (.A1(_15149_),
    .A2(_02494_),
    .A3(_02496_),
    .ZN(_02497_));
 OAI21_X1 _25481_ (.A(_02486_),
    .B1(_02493_),
    .B2(_02497_),
    .ZN(_02498_));
 NAND2_X1 _25482_ (.A1(_02296_),
    .A2(_02343_),
    .ZN(_02499_));
 AOI21_X1 _25483_ (.A(_02426_),
    .B1(_02415_),
    .B2(_02390_),
    .ZN(_02500_));
 AND2_X1 _25484_ (.A1(_02499_),
    .A2(_02500_),
    .ZN(_02501_));
 NOR3_X1 _25485_ (.A1(_15142_),
    .A2(_02450_),
    .A3(_02454_),
    .ZN(_02502_));
 OAI21_X1 _25486_ (.A(_02449_),
    .B1(_02501_),
    .B2(_02502_),
    .ZN(_02503_));
 XNOR2_X2 _25487_ (.A(_06567_),
    .B(_02329_),
    .ZN(_02504_));
 NAND2_X1 _25488_ (.A1(_02447_),
    .A2(_02504_),
    .ZN(_02505_));
 NAND2_X4 _25489_ (.A1(_02296_),
    .A2(net1095),
    .ZN(_02506_));
 OAI21_X1 _25490_ (.A(_02506_),
    .B1(_15133_),
    .B2(net1044),
    .ZN(_02507_));
 XNOR2_X1 _25491_ (.A(_02440_),
    .B(_02507_),
    .ZN(_02508_));
 CLKBUF_X3 _25492_ (.A(_02362_),
    .Z(_02509_));
 NOR2_X1 _25493_ (.A1(_02396_),
    .A2(_02509_),
    .ZN(_02510_));
 AOI21_X1 _25494_ (.A(_02505_),
    .B1(_02508_),
    .B2(_02510_),
    .ZN(_02511_));
 NAND4_X2 _25495_ (.A1(_02492_),
    .A2(_02498_),
    .A3(_02503_),
    .A4(_02511_),
    .ZN(_02512_));
 NAND4_X4 _25496_ (.A1(_02410_),
    .A2(_02488_),
    .A3(_02446_),
    .A4(_02512_),
    .ZN(_00112_));
 NAND2_X1 _25497_ (.A1(_02399_),
    .A2(_02391_),
    .ZN(_02513_));
 NAND3_X1 _25498_ (.A1(_02426_),
    .A2(_02499_),
    .A3(_02513_),
    .ZN(_02514_));
 NOR2_X1 _25499_ (.A1(_02406_),
    .A2(_02311_),
    .ZN(_02515_));
 AOI221_X2 _25500_ (.A(_02361_),
    .B1(_02403_),
    .B2(_02515_),
    .C1(_02483_),
    .C2(net143),
    .ZN(_02516_));
 AOI221_X2 _25501_ (.A(_02419_),
    .B1(_02484_),
    .B2(_02295_),
    .C1(_02386_),
    .C2(net144),
    .ZN(_02517_));
 BUF_X4 _25502_ (.A(_02361_),
    .Z(_02518_));
 BUF_X4 _25503_ (.A(_02518_),
    .Z(_02519_));
 AOI221_X1 _25504_ (.A(_02447_),
    .B1(_02514_),
    .B2(_02516_),
    .C1(_02517_),
    .C2(_02519_),
    .ZN(_02520_));
 INV_X4 _25505_ (.A(net588),
    .ZN(_02521_));
 NAND2_X2 _25506_ (.A1(_02521_),
    .A2(_02379_),
    .ZN(_02522_));
 NAND2_X1 _25507_ (.A1(_02399_),
    .A2(_02403_),
    .ZN(_02523_));
 AOI21_X1 _25508_ (.A(_02427_),
    .B1(_02522_),
    .B2(_02523_),
    .ZN(_02524_));
 NAND2_X1 _25509_ (.A1(_02509_),
    .A2(_02325_),
    .ZN(_02525_));
 NAND2_X2 _25510_ (.A1(_02311_),
    .A2(_02349_),
    .ZN(_02526_));
 NOR2_X1 _25511_ (.A1(_02443_),
    .A2(_02526_),
    .ZN(_02527_));
 NAND2_X1 _25512_ (.A1(net1040),
    .A2(_02350_),
    .ZN(_02528_));
 AOI21_X1 _25513_ (.A(_02313_),
    .B1(_02496_),
    .B2(_02528_),
    .ZN(_02529_));
 NAND2_X1 _25514_ (.A1(_02384_),
    .A2(_02447_),
    .ZN(_02530_));
 NAND2_X1 _25515_ (.A1(net580),
    .A2(_02426_),
    .ZN(_02531_));
 NOR2_X1 _25516_ (.A1(_02440_),
    .A2(_02531_),
    .ZN(_02532_));
 OAI33_X1 _25517_ (.A1(_02524_),
    .A2(_02525_),
    .A3(_02527_),
    .B1(_02529_),
    .B2(_02530_),
    .B3(_02532_),
    .ZN(_02533_));
 OR3_X2 _25518_ (.A1(_02414_),
    .A2(_02520_),
    .A3(_02533_),
    .ZN(_02534_));
 NAND2_X1 _25519_ (.A1(_02369_),
    .A2(_02433_),
    .ZN(_02535_));
 NAND2_X2 _25520_ (.A1(net731),
    .A2(_02317_),
    .ZN(_02536_));
 NOR2_X2 _25521_ (.A1(net590),
    .A2(_02316_),
    .ZN(_02537_));
 NOR2_X1 _25522_ (.A1(_02415_),
    .A2(_02537_),
    .ZN(_02538_));
 INV_X1 _25523_ (.A(_15154_),
    .ZN(_02539_));
 AOI221_X2 _25524_ (.A(_02535_),
    .B1(_02536_),
    .B2(_02538_),
    .C1(_02416_),
    .C2(_02539_),
    .ZN(_02540_));
 NAND2_X1 _25525_ (.A1(_02422_),
    .A2(_02440_),
    .ZN(_02541_));
 AOI21_X2 _25526_ (.A(_02402_),
    .B1(_02350_),
    .B2(_02521_),
    .ZN(_02542_));
 AOI21_X1 _25527_ (.A(_02530_),
    .B1(_02541_),
    .B2(_02542_),
    .ZN(_02543_));
 NOR2_X4 _25528_ (.A1(_02296_),
    .A2(net1174),
    .ZN(_02544_));
 OAI21_X1 _25529_ (.A(_15149_),
    .B1(_02386_),
    .B2(_02544_),
    .ZN(_02545_));
 AOI21_X1 _25530_ (.A(_02540_),
    .B1(_02543_),
    .B2(_02545_),
    .ZN(_02546_));
 NAND2_X4 _25531_ (.A1(_02361_),
    .A2(_02433_),
    .ZN(_02547_));
 CLKBUF_X3 _25532_ (.A(_02316_),
    .Z(_02548_));
 NAND2_X1 _25533_ (.A1(net580),
    .A2(_02548_),
    .ZN(_02549_));
 AOI21_X1 _25534_ (.A(_02376_),
    .B1(_02418_),
    .B2(_02549_),
    .ZN(_02550_));
 NOR2_X1 _25535_ (.A1(_02547_),
    .A2(_02550_),
    .ZN(_02551_));
 NOR2_X2 _25536_ (.A1(_02346_),
    .A2(_02344_),
    .ZN(_02552_));
 OAI21_X1 _25537_ (.A(_02427_),
    .B1(_02552_),
    .B2(_02455_),
    .ZN(_02553_));
 NOR2_X2 _25538_ (.A1(_02295_),
    .A2(_02391_),
    .ZN(_02554_));
 AOI21_X1 _25539_ (.A(_02525_),
    .B1(_02554_),
    .B2(net145),
    .ZN(_02555_));
 AOI221_X2 _25540_ (.A(_02396_),
    .B1(_02424_),
    .B2(_02551_),
    .C1(_02553_),
    .C2(_02555_),
    .ZN(_02556_));
 AOI21_X2 _25541_ (.A(_02504_),
    .B1(_02546_),
    .B2(_02556_),
    .ZN(_02557_));
 OAI221_X2 _25542_ (.A(_02383_),
    .B1(_02404_),
    .B2(_02296_),
    .C1(_02522_),
    .C2(_02318_),
    .ZN(_02558_));
 NAND2_X1 _25543_ (.A1(_02405_),
    .A2(_02379_),
    .ZN(_02559_));
 AOI21_X1 _25544_ (.A(_02427_),
    .B1(_02345_),
    .B2(_02559_),
    .ZN(_02560_));
 OAI21_X1 _25545_ (.A(_02319_),
    .B1(_02440_),
    .B2(_02422_),
    .ZN(_02561_));
 OAI21_X1 _25546_ (.A(_02313_),
    .B1(_02400_),
    .B2(_02405_),
    .ZN(_02562_));
 NOR2_X4 _25547_ (.A1(net720),
    .A2(_02342_),
    .ZN(_02563_));
 OAI22_X1 _25548_ (.A1(_02544_),
    .A2(_02561_),
    .B1(_02562_),
    .B2(_02563_),
    .ZN(_02564_));
 OAI221_X1 _25549_ (.A(_02447_),
    .B1(_02558_),
    .B2(_02560_),
    .C1(_02564_),
    .C2(_02384_),
    .ZN(_02565_));
 NAND2_X1 _25550_ (.A1(_02442_),
    .A2(_02350_),
    .ZN(_02566_));
 AOI21_X1 _25551_ (.A(_02548_),
    .B1(_02376_),
    .B2(_02332_),
    .ZN(_02567_));
 NAND2_X1 _25552_ (.A1(_02453_),
    .A2(_02403_),
    .ZN(_02568_));
 AOI221_X1 _25553_ (.A(_02509_),
    .B1(_02566_),
    .B2(_02567_),
    .C1(_02568_),
    .C2(_02500_),
    .ZN(_02569_));
 NAND2_X1 _25554_ (.A1(_02442_),
    .A2(_02375_),
    .ZN(_02570_));
 AOI221_X2 _25555_ (.A(_02475_),
    .B1(_02542_),
    .B2(_02570_),
    .C1(_02490_),
    .C2(_02313_),
    .ZN(_02571_));
 OAI21_X1 _25556_ (.A(_02435_),
    .B1(_02569_),
    .B2(_02571_),
    .ZN(_02572_));
 NAND3_X1 _25557_ (.A1(_02397_),
    .A2(_02565_),
    .A3(_02572_),
    .ZN(_02573_));
 OAI21_X1 _25558_ (.A(_02519_),
    .B1(_02440_),
    .B2(_15150_),
    .ZN(_02574_));
 NAND2_X1 _25559_ (.A1(_02435_),
    .A2(_02574_),
    .ZN(_02575_));
 MUX2_X2 _25560_ (.A(_02371_),
    .B(_02442_),
    .S(_02317_),
    .Z(_02576_));
 NAND2_X2 _25561_ (.A1(_02362_),
    .A2(_02343_),
    .ZN(_02577_));
 NAND3_X1 _25562_ (.A1(_02443_),
    .A2(_02319_),
    .A3(_02400_),
    .ZN(_02578_));
 NAND2_X4 _25563_ (.A1(_02316_),
    .A2(_02403_),
    .ZN(_02579_));
 OAI221_X2 _25564_ (.A(_02578_),
    .B1(_02562_),
    .B2(_02552_),
    .C1(_15133_),
    .C2(_02579_),
    .ZN(_02580_));
 OAI221_X2 _25565_ (.A(_02575_),
    .B1(_02576_),
    .B2(_02577_),
    .C1(_02580_),
    .C2(_02519_),
    .ZN(_02581_));
 NOR2_X4 _25566_ (.A1(_02362_),
    .A2(_02325_),
    .ZN(_02582_));
 XNOR2_X2 _25567_ (.A(_02314_),
    .B(_02403_),
    .ZN(_02583_));
 OAI22_X1 _25568_ (.A1(_02544_),
    .A2(_02561_),
    .B1(_02583_),
    .B2(_15142_),
    .ZN(_02584_));
 AOI21_X1 _25569_ (.A(_02397_),
    .B1(_02582_),
    .B2(_02584_),
    .ZN(_02585_));
 AOI21_X2 _25570_ (.A(_02436_),
    .B1(_02581_),
    .B2(_02585_),
    .ZN(_02586_));
 AOI22_X4 _25571_ (.A1(_02534_),
    .A2(_02557_),
    .B1(_02573_),
    .B2(_02586_),
    .ZN(_00113_));
 NAND2_X2 _25572_ (.A1(_02356_),
    .A2(_02504_),
    .ZN(_02587_));
 INV_X1 _25573_ (.A(_02587_),
    .ZN(_02588_));
 NAND2_X1 _25574_ (.A1(net732),
    .A2(_02375_),
    .ZN(_02589_));
 AOI21_X1 _25575_ (.A(_02548_),
    .B1(_02589_),
    .B2(_02566_),
    .ZN(_02590_));
 NOR2_X4 _25576_ (.A1(_02369_),
    .A2(_02433_),
    .ZN(_02591_));
 OAI21_X1 _25577_ (.A(_02591_),
    .B1(_02444_),
    .B2(net1042),
    .ZN(_02592_));
 AOI21_X1 _25578_ (.A(_02350_),
    .B1(_02316_),
    .B2(net1040),
    .ZN(_02593_));
 AND2_X1 _25579_ (.A1(_02418_),
    .A2(_02593_),
    .ZN(_02594_));
 AOI21_X4 _25580_ (.A(_02383_),
    .B1(net719),
    .B2(_02379_),
    .ZN(_02595_));
 NAND2_X2 _25581_ (.A1(_02595_),
    .A2(_02434_),
    .ZN(_02596_));
 OAI221_X2 _25582_ (.A(_02588_),
    .B1(_02590_),
    .B2(_02592_),
    .C1(_02596_),
    .C2(_02594_),
    .ZN(_02597_));
 BUF_X4 _25583_ (.A(_02402_),
    .Z(_02598_));
 NOR3_X2 _25584_ (.A1(_02598_),
    .A2(_02386_),
    .A3(_02471_),
    .ZN(_02599_));
 NOR2_X1 _25585_ (.A1(_02332_),
    .A2(_02375_),
    .ZN(_02600_));
 NOR3_X1 _25586_ (.A1(_02318_),
    .A2(_02385_),
    .A3(_02600_),
    .ZN(_02601_));
 NOR2_X2 _25587_ (.A1(_02601_),
    .A2(_02599_),
    .ZN(_02602_));
 NOR2_X4 _25588_ (.A1(_02361_),
    .A2(_02433_),
    .ZN(_02603_));
 AND2_X1 _25589_ (.A1(_02351_),
    .A2(_02568_),
    .ZN(_02604_));
 NOR2_X2 _25590_ (.A1(net590),
    .A2(_02349_),
    .ZN(_02605_));
 NOR2_X1 _25591_ (.A1(_02563_),
    .A2(_02605_),
    .ZN(_02606_));
 MUX2_X1 _25592_ (.A(_02604_),
    .B(_02606_),
    .S(_02318_),
    .Z(_02607_));
 AOI221_X2 _25593_ (.A(_02597_),
    .B1(_02603_),
    .B2(_02602_),
    .C1(_02607_),
    .C2(_02582_),
    .ZN(_02608_));
 NAND2_X1 _25594_ (.A1(_02332_),
    .A2(_02422_),
    .ZN(_02609_));
 AOI221_X1 _25595_ (.A(_02372_),
    .B1(_02483_),
    .B2(_02609_),
    .C1(_02484_),
    .C2(_02495_),
    .ZN(_02610_));
 MUX2_X1 _25596_ (.A(net143),
    .B(_02406_),
    .S(_02342_),
    .Z(_02611_));
 AOI22_X1 _25597_ (.A1(_02399_),
    .A2(_02364_),
    .B1(_02611_),
    .B2(_02548_),
    .ZN(_02612_));
 MUX2_X1 _25598_ (.A(_02610_),
    .B(_02612_),
    .S(_02518_),
    .Z(_02613_));
 NAND2_X1 _25599_ (.A1(_02346_),
    .A2(_02312_),
    .ZN(_02614_));
 AND3_X1 _25600_ (.A1(_02383_),
    .A2(_02614_),
    .A3(_02536_),
    .ZN(_02615_));
 OAI21_X1 _25601_ (.A(_02415_),
    .B1(_02475_),
    .B2(_15145_),
    .ZN(_02616_));
 MUX2_X1 _25602_ (.A(_15156_),
    .B(_02614_),
    .S(_02362_),
    .Z(_02617_));
 OAI22_X1 _25603_ (.A1(_02615_),
    .A2(_02616_),
    .B1(_02617_),
    .B2(_02400_),
    .ZN(_02618_));
 MUX2_X1 _25604_ (.A(_02613_),
    .B(_02618_),
    .S(_02435_),
    .Z(_02619_));
 NOR2_X1 _25605_ (.A1(_02396_),
    .A2(_02504_),
    .ZN(_02620_));
 NAND2_X2 _25606_ (.A1(_02395_),
    .A2(_02361_),
    .ZN(_02621_));
 NOR2_X1 _25607_ (.A1(_02435_),
    .A2(_02621_),
    .ZN(_02622_));
 OAI21_X1 _25608_ (.A(_02318_),
    .B1(_02376_),
    .B2(_02390_),
    .ZN(_02623_));
 NOR2_X1 _25609_ (.A1(_02521_),
    .A2(_02376_),
    .ZN(_02624_));
 OAI21_X1 _25610_ (.A(_02426_),
    .B1(_02380_),
    .B2(_02366_),
    .ZN(_02625_));
 OAI221_X2 _25611_ (.A(_02622_),
    .B1(_02623_),
    .B2(_02544_),
    .C1(_02624_),
    .C2(_02625_),
    .ZN(_02626_));
 NAND2_X1 _25612_ (.A1(_02366_),
    .A2(_02316_),
    .ZN(_02627_));
 AOI21_X1 _25613_ (.A(_02400_),
    .B1(_02531_),
    .B2(_02627_),
    .ZN(_02628_));
 NAND2_X1 _25614_ (.A1(net590),
    .A2(_02311_),
    .ZN(_02629_));
 AOI21_X1 _25615_ (.A(_02411_),
    .B1(_02506_),
    .B2(_02629_),
    .ZN(_02630_));
 OAI21_X1 _25616_ (.A(_02384_),
    .B1(_02628_),
    .B2(_02630_),
    .ZN(_02631_));
 NOR2_X1 _25617_ (.A1(_02475_),
    .A2(_02537_),
    .ZN(_02632_));
 MUX2_X1 _25618_ (.A(_02366_),
    .B(net1044),
    .S(_02380_),
    .Z(_02633_));
 OAI21_X1 _25619_ (.A(_02632_),
    .B1(_02633_),
    .B2(_02427_),
    .ZN(_02634_));
 NAND4_X1 _25620_ (.A1(_02397_),
    .A2(_02435_),
    .A3(_02631_),
    .A4(_02634_),
    .ZN(_02635_));
 BUF_X4 _25621_ (.A(_02317_),
    .Z(_02636_));
 NAND2_X1 _25622_ (.A1(_15136_),
    .A2(_02461_),
    .ZN(_02637_));
 NAND2_X1 _25623_ (.A1(_15136_),
    .A2(_02459_),
    .ZN(_02638_));
 MUX2_X2 _25624_ (.A(_02637_),
    .B(_02638_),
    .S(_02339_),
    .Z(_02639_));
 INV_X4 _25625_ (.A(_15136_),
    .ZN(_02640_));
 NOR3_X2 _25626_ (.A1(_02333_),
    .A2(_02640_),
    .A3(_02467_),
    .ZN(_02641_));
 NOR3_X2 _25627_ (.A1(_02464_),
    .A2(_02640_),
    .A3(_02466_),
    .ZN(_02642_));
 NOR2_X2 _25628_ (.A1(_02641_),
    .A2(_02642_),
    .ZN(_02643_));
 NAND3_X1 _25629_ (.A1(_02636_),
    .A2(_02639_),
    .A3(_02643_),
    .ZN(_02644_));
 OAI21_X1 _25630_ (.A(_02313_),
    .B1(_02400_),
    .B2(_02453_),
    .ZN(_02645_));
 NOR2_X1 _25631_ (.A1(_02279_),
    .A2(_02375_),
    .ZN(_02646_));
 OAI22_X1 _25632_ (.A1(_02554_),
    .A2(_02644_),
    .B1(_02645_),
    .B2(_02646_),
    .ZN(_02647_));
 AOI21_X1 _25633_ (.A(_02436_),
    .B1(_02603_),
    .B2(_02647_),
    .ZN(_02648_));
 OAI211_X2 _25634_ (.A(_02626_),
    .B(_02635_),
    .C1(_02648_),
    .C2(_02414_),
    .ZN(_02649_));
 NAND3_X1 _25635_ (.A1(net144),
    .A2(_02295_),
    .A3(_02434_),
    .ZN(_02650_));
 NAND2_X1 _25636_ (.A1(_02380_),
    .A2(_02650_),
    .ZN(_02651_));
 MUX2_X1 _25637_ (.A(_02346_),
    .B(net1040),
    .S(_02433_),
    .Z(_02652_));
 AOI221_X2 _25638_ (.A(_02651_),
    .B1(_02472_),
    .B2(_02325_),
    .C1(_02636_),
    .C2(_02652_),
    .ZN(_02653_));
 NAND2_X1 _25639_ (.A1(_15150_),
    .A2(_02434_),
    .ZN(_02654_));
 OAI21_X1 _25640_ (.A(_02654_),
    .B1(_02434_),
    .B2(_15147_),
    .ZN(_02655_));
 OAI21_X1 _25641_ (.A(_02519_),
    .B1(_02416_),
    .B2(_02655_),
    .ZN(_02656_));
 NAND3_X1 _25642_ (.A1(net145),
    .A2(_02400_),
    .A3(_02506_),
    .ZN(_02657_));
 MUX2_X1 _25643_ (.A(_02548_),
    .B(_02380_),
    .S(net1040),
    .Z(_02658_));
 OAI221_X2 _25644_ (.A(_02657_),
    .B1(_02536_),
    .B2(_02386_),
    .C1(_02521_),
    .C2(_02658_),
    .ZN(_02659_));
 NOR3_X1 _25645_ (.A1(_02427_),
    .A2(_02388_),
    .A3(_02455_),
    .ZN(_02660_));
 OAI21_X1 _25646_ (.A(_02434_),
    .B1(_02611_),
    .B2(_02319_),
    .ZN(_02661_));
 OAI22_X2 _25647_ (.A1(_02435_),
    .A2(_02659_),
    .B1(_02660_),
    .B2(_02661_),
    .ZN(_02662_));
 OAI221_X2 _25648_ (.A(_02436_),
    .B1(_02653_),
    .B2(_02656_),
    .C1(_02662_),
    .C2(_02519_),
    .ZN(_02663_));
 AOI221_X2 _25649_ (.A(_02608_),
    .B1(_02619_),
    .B2(_02620_),
    .C1(_02649_),
    .C2(_02663_),
    .ZN(_00114_));
 OAI21_X1 _25650_ (.A(_02427_),
    .B1(_02454_),
    .B2(_02554_),
    .ZN(_02664_));
 AOI21_X2 _25651_ (.A(_02311_),
    .B1(_02341_),
    .B2(_02521_),
    .ZN(_02665_));
 NOR2_X2 _25652_ (.A1(_02378_),
    .A2(net718),
    .ZN(_02666_));
 NAND2_X1 _25653_ (.A1(_02379_),
    .A2(_02666_),
    .ZN(_02667_));
 AOI21_X1 _25654_ (.A(_02547_),
    .B1(_02665_),
    .B2(_02667_),
    .ZN(_02668_));
 NOR2_X2 _25655_ (.A1(_02380_),
    .A2(_02506_),
    .ZN(_02669_));
 XNOR2_X1 _25656_ (.A(_02426_),
    .B(_02376_),
    .ZN(_02670_));
 AOI21_X1 _25657_ (.A(_02669_),
    .B1(_02670_),
    .B2(_02366_),
    .ZN(_02671_));
 AOI22_X1 _25658_ (.A1(_02664_),
    .A2(_02668_),
    .B1(_02671_),
    .B2(_02591_),
    .ZN(_02672_));
 AOI21_X1 _25659_ (.A(_02324_),
    .B1(_02312_),
    .B2(_02371_),
    .ZN(_02673_));
 AOI221_X2 _25660_ (.A(_02518_),
    .B1(_02593_),
    .B2(_02673_),
    .C1(_02483_),
    .C2(_02378_),
    .ZN(_02674_));
 MUX2_X1 _25661_ (.A(_02526_),
    .B(_02579_),
    .S(_02325_),
    .Z(_02675_));
 OAI21_X1 _25662_ (.A(_02674_),
    .B1(_02675_),
    .B2(_02390_),
    .ZN(_02676_));
 AOI21_X1 _25663_ (.A(_02587_),
    .B1(_02672_),
    .B2(_02676_),
    .ZN(_02677_));
 NAND2_X1 _25664_ (.A1(net143),
    .A2(_02349_),
    .ZN(_02678_));
 NOR2_X1 _25665_ (.A1(_02316_),
    .A2(_02544_),
    .ZN(_02679_));
 AOI21_X1 _25666_ (.A(_02312_),
    .B1(_02375_),
    .B2(_02371_),
    .ZN(_02680_));
 AOI221_X2 _25667_ (.A(_02362_),
    .B1(_02678_),
    .B2(_02679_),
    .C1(_02680_),
    .C2(_02559_),
    .ZN(_02681_));
 NAND3_X1 _25668_ (.A1(_02426_),
    .A2(_02518_),
    .A3(_02513_),
    .ZN(_02682_));
 NOR2_X1 _25669_ (.A1(_02455_),
    .A2(_02682_),
    .ZN(_02683_));
 NAND2_X1 _25670_ (.A1(_02318_),
    .A2(_02518_),
    .ZN(_02684_));
 NOR3_X1 _25671_ (.A1(_02392_),
    .A2(_02454_),
    .A3(_02684_),
    .ZN(_02685_));
 OR4_X1 _25672_ (.A1(_02435_),
    .A2(_02681_),
    .A3(_02683_),
    .A4(_02685_),
    .ZN(_02686_));
 AOI21_X1 _25673_ (.A(_02319_),
    .B1(_02473_),
    .B2(_02522_),
    .ZN(_02687_));
 OAI21_X1 _25674_ (.A(_02582_),
    .B1(_02579_),
    .B2(_15133_),
    .ZN(_02688_));
 OAI21_X1 _25675_ (.A(_02620_),
    .B1(_02687_),
    .B2(_02688_),
    .ZN(_02689_));
 NOR2_X2 _25676_ (.A1(net720),
    .A2(_02548_),
    .ZN(_02690_));
 AOI22_X1 _25677_ (.A1(_02690_),
    .A2(_02490_),
    .B1(_02506_),
    .B2(_02385_),
    .ZN(_02691_));
 NAND2_X1 _25678_ (.A1(_02390_),
    .A2(_02483_),
    .ZN(_02692_));
 AOI21_X1 _25679_ (.A(_02547_),
    .B1(_02691_),
    .B2(_02692_),
    .ZN(_02693_));
 NOR2_X1 _25680_ (.A1(_02689_),
    .A2(_02693_),
    .ZN(_02694_));
 OAI21_X1 _25681_ (.A(_02506_),
    .B1(_02296_),
    .B2(net144),
    .ZN(_02695_));
 AOI221_X2 _25682_ (.A(_02547_),
    .B1(_02695_),
    .B2(_02341_),
    .C1(_02364_),
    .C2(net732),
    .ZN(_02696_));
 AOI21_X1 _25683_ (.A(_02324_),
    .B1(_02348_),
    .B2(_02279_),
    .ZN(_02697_));
 AOI21_X1 _25684_ (.A(_02324_),
    .B1(_02341_),
    .B2(_02366_),
    .ZN(_02698_));
 AOI21_X2 _25685_ (.A(_02315_),
    .B1(net1175),
    .B2(net1042),
    .ZN(_02699_));
 AOI221_X2 _25686_ (.A(_02361_),
    .B1(_02665_),
    .B2(_02697_),
    .C1(_02698_),
    .C2(_02699_),
    .ZN(_02700_));
 NOR2_X1 _25687_ (.A1(net143),
    .A2(_02311_),
    .ZN(_02701_));
 AOI21_X1 _25688_ (.A(_02433_),
    .B1(_02701_),
    .B2(_02403_),
    .ZN(_02702_));
 MUX2_X1 _25689_ (.A(_02371_),
    .B(_02295_),
    .S(_02348_),
    .Z(_02703_));
 OAI221_X2 _25690_ (.A(_02702_),
    .B1(_02703_),
    .B2(_02316_),
    .C1(_02528_),
    .C2(_02296_),
    .ZN(_02704_));
 MUX2_X1 _25691_ (.A(_02371_),
    .B(_02442_),
    .S(_02342_),
    .Z(_02705_));
 OAI21_X2 _25692_ (.A(_02402_),
    .B1(_02350_),
    .B2(net143),
    .ZN(_02706_));
 NOR2_X2 _25693_ (.A1(_02374_),
    .A2(_02342_),
    .ZN(_02707_));
 OAI22_X2 _25694_ (.A1(_02598_),
    .A2(_02705_),
    .B1(_02706_),
    .B2(_02707_),
    .ZN(_02708_));
 AOI221_X2 _25695_ (.A(_02696_),
    .B1(_02700_),
    .B2(_02704_),
    .C1(_02708_),
    .C2(_02591_),
    .ZN(_02709_));
 NOR3_X1 _25696_ (.A1(_15133_),
    .A2(_02391_),
    .A3(_02325_),
    .ZN(_02710_));
 NAND4_X4 _25697_ (.A1(_02470_),
    .A2(_02463_),
    .A3(_02639_),
    .A4(net1097),
    .ZN(_02711_));
 OAI21_X4 _25698_ (.A(_02548_),
    .B1(_02711_),
    .B2(_02434_),
    .ZN(_02712_));
 OAI21_X1 _25699_ (.A(_02426_),
    .B1(_02380_),
    .B2(net1043),
    .ZN(_02713_));
 NOR3_X1 _25700_ (.A1(_15122_),
    .A2(_02376_),
    .A3(_02434_),
    .ZN(_02714_));
 OAI221_X2 _25701_ (.A(_02475_),
    .B1(_02712_),
    .B2(_02710_),
    .C1(_02713_),
    .C2(_02714_),
    .ZN(_02715_));
 OAI221_X1 _25702_ (.A(_02591_),
    .B1(_02404_),
    .B2(net145),
    .C1(_02405_),
    .C2(_02444_),
    .ZN(_02716_));
 AOI21_X1 _25703_ (.A(_15122_),
    .B1(_02636_),
    .B2(_02473_),
    .ZN(_02717_));
 NOR2_X1 _25704_ (.A1(_02598_),
    .A2(_02666_),
    .ZN(_02718_));
 NOR2_X4 _25705_ (.A1(_02640_),
    .A2(net1096),
    .ZN(_02719_));
 OAI21_X1 _25706_ (.A(_02415_),
    .B1(_02718_),
    .B2(_02719_),
    .ZN(_02720_));
 OAI21_X1 _25707_ (.A(_02720_),
    .B1(_02576_),
    .B2(_02400_),
    .ZN(_02721_));
 OAI221_X1 _25708_ (.A(_02715_),
    .B1(_02716_),
    .B2(_02717_),
    .C1(_02721_),
    .C2(_02547_),
    .ZN(_02722_));
 MUX2_X1 _25709_ (.A(_02709_),
    .B(_02722_),
    .S(_02504_),
    .Z(_02723_));
 AOI221_X2 _25710_ (.A(_02677_),
    .B1(_02686_),
    .B2(_02694_),
    .C1(_02723_),
    .C2(_02397_),
    .ZN(_00115_));
 OAI221_X2 _25711_ (.A(_02427_),
    .B1(_02519_),
    .B2(_02583_),
    .C1(_02577_),
    .C2(net581),
    .ZN(_02724_));
 NOR2_X1 _25712_ (.A1(_02509_),
    .A2(_02411_),
    .ZN(_02725_));
 MUX2_X1 _25713_ (.A(_02407_),
    .B(_15122_),
    .S(_02518_),
    .Z(_02726_));
 AOI22_X1 _25714_ (.A1(_02399_),
    .A2(_02725_),
    .B1(_02726_),
    .B2(_02440_),
    .ZN(_02727_));
 OAI211_X2 _25715_ (.A(_02397_),
    .B(_02724_),
    .C1(_02727_),
    .C2(_15149_),
    .ZN(_02728_));
 NAND2_X2 _25716_ (.A1(_02643_),
    .A2(_02639_),
    .ZN(_02729_));
 NOR2_X1 _25717_ (.A1(_02407_),
    .A2(_02548_),
    .ZN(_02730_));
 NOR4_X1 _25718_ (.A1(_02475_),
    .A2(_02415_),
    .A3(_02477_),
    .A4(_02730_),
    .ZN(_02731_));
 NAND2_X1 _25719_ (.A1(net1044),
    .A2(_02356_),
    .ZN(_02732_));
 OAI33_X1 _25720_ (.A1(_15142_),
    .A2(_02370_),
    .A3(_02729_),
    .B1(_02725_),
    .B2(_02731_),
    .B3(_02732_),
    .ZN(_02733_));
 NAND2_X1 _25721_ (.A1(_15122_),
    .A2(_02733_),
    .ZN(_02734_));
 OAI21_X1 _25722_ (.A(_02414_),
    .B1(_02477_),
    .B2(_02730_),
    .ZN(_02735_));
 NOR2_X1 _25723_ (.A1(_02577_),
    .A2(_02735_),
    .ZN(_02736_));
 NOR3_X1 _25724_ (.A1(_02370_),
    .A2(_02458_),
    .A3(_02729_),
    .ZN(_02737_));
 NOR3_X1 _25725_ (.A1(_02447_),
    .A2(_02736_),
    .A3(_02737_),
    .ZN(_02738_));
 AOI22_X1 _25726_ (.A1(_02319_),
    .A2(_02519_),
    .B1(_02440_),
    .B2(_02407_),
    .ZN(_02739_));
 OAI21_X1 _25727_ (.A(_02384_),
    .B1(_02440_),
    .B2(_02719_),
    .ZN(_02740_));
 NAND4_X1 _25728_ (.A1(_15133_),
    .A2(_02414_),
    .A3(_02739_),
    .A4(_02740_),
    .ZN(_02741_));
 NAND4_X1 _25729_ (.A1(_02728_),
    .A2(_02734_),
    .A3(_02738_),
    .A4(_02741_),
    .ZN(_02742_));
 OAI221_X1 _25730_ (.A(_02578_),
    .B1(_02706_),
    .B2(_02386_),
    .C1(_02579_),
    .C2(_02399_),
    .ZN(_02743_));
 NOR2_X1 _25731_ (.A1(_02521_),
    .A2(_02636_),
    .ZN(_02744_));
 NAND2_X1 _25732_ (.A1(_02416_),
    .A2(_02744_),
    .ZN(_02745_));
 AOI21_X1 _25733_ (.A(_02396_),
    .B1(_02440_),
    .B2(_02443_),
    .ZN(_02746_));
 AOI21_X1 _25734_ (.A(_02384_),
    .B1(_02745_),
    .B2(_02746_),
    .ZN(_02747_));
 NAND2_X1 _25735_ (.A1(_02427_),
    .A2(_02396_),
    .ZN(_02748_));
 AOI21_X1 _25736_ (.A(_02748_),
    .B1(_02566_),
    .B2(_02345_),
    .ZN(_02749_));
 OAI22_X1 _25737_ (.A1(_02621_),
    .A2(_02743_),
    .B1(_02747_),
    .B2(_02749_),
    .ZN(_02750_));
 OAI21_X1 _25738_ (.A(_15142_),
    .B1(_02450_),
    .B2(_02563_),
    .ZN(_02751_));
 AOI21_X1 _25739_ (.A(_02370_),
    .B1(_02364_),
    .B2(_02366_),
    .ZN(_02752_));
 AOI21_X1 _25740_ (.A(_02435_),
    .B1(_02751_),
    .B2(_02752_),
    .ZN(_02753_));
 AOI21_X1 _25741_ (.A(_02436_),
    .B1(_02750_),
    .B2(_02753_),
    .ZN(_02754_));
 MUX2_X1 _25742_ (.A(_02453_),
    .B(net144),
    .S(_02349_),
    .Z(_02755_));
 NOR2_X1 _25743_ (.A1(_02319_),
    .A2(_02755_),
    .ZN(_02756_));
 NOR3_X1 _25744_ (.A1(_02313_),
    .A2(_02707_),
    .A3(_02605_),
    .ZN(_02757_));
 OR3_X1 _25745_ (.A1(_02519_),
    .A2(_02756_),
    .A3(_02757_),
    .ZN(_02758_));
 OAI21_X1 _25746_ (.A(_02416_),
    .B1(_02428_),
    .B2(_02690_),
    .ZN(_02759_));
 NAND3_X2 _25747_ (.A1(_02519_),
    .A2(_02424_),
    .A3(_02759_),
    .ZN(_02760_));
 NAND3_X2 _25748_ (.A1(_02414_),
    .A2(_02758_),
    .A3(_02760_),
    .ZN(_02761_));
 NAND2_X1 _25749_ (.A1(_02295_),
    .A2(_02379_),
    .ZN(_02762_));
 NOR2_X1 _25750_ (.A1(net1044),
    .A2(_02762_),
    .ZN(_02763_));
 OAI21_X1 _25751_ (.A(_02439_),
    .B1(_02484_),
    .B2(net145),
    .ZN(_02764_));
 NOR3_X1 _25752_ (.A1(_02669_),
    .A2(_02763_),
    .A3(_02764_),
    .ZN(_02765_));
 NAND2_X1 _25753_ (.A1(_02314_),
    .A2(_02316_),
    .ZN(_02766_));
 NAND2_X1 _25754_ (.A1(_02449_),
    .A2(_02766_),
    .ZN(_02767_));
 AOI221_X2 _25755_ (.A(_02767_),
    .B1(_02554_),
    .B2(net1044),
    .C1(_02405_),
    .C2(_02364_),
    .ZN(_02768_));
 NOR3_X2 _25756_ (.A1(_02437_),
    .A2(_02765_),
    .A3(_02768_),
    .ZN(_02769_));
 NOR2_X1 _25757_ (.A1(_02407_),
    .A2(_02416_),
    .ZN(_02770_));
 NOR3_X1 _25758_ (.A1(_02319_),
    .A2(_02770_),
    .A3(_02563_),
    .ZN(_02771_));
 NAND2_X1 _25759_ (.A1(_02397_),
    .A2(_02506_),
    .ZN(_02772_));
 MUX2_X1 _25760_ (.A(_02604_),
    .B(_02711_),
    .S(_02427_),
    .Z(_02773_));
 OAI221_X2 _25761_ (.A(_02519_),
    .B1(_02771_),
    .B2(_02772_),
    .C1(_02773_),
    .C2(_02397_),
    .ZN(_02774_));
 XNOR2_X1 _25762_ (.A(_02426_),
    .B(_02356_),
    .ZN(_02775_));
 OAI221_X1 _25763_ (.A(_02384_),
    .B1(_02345_),
    .B2(_02414_),
    .C1(_02775_),
    .C2(_02366_),
    .ZN(_02776_));
 OAI21_X1 _25764_ (.A(_02411_),
    .B1(_02396_),
    .B2(_02422_),
    .ZN(_02777_));
 OAI21_X1 _25765_ (.A(_02777_),
    .B1(_02522_),
    .B2(_02396_),
    .ZN(_02778_));
 AOI21_X1 _25766_ (.A(_02776_),
    .B1(_02778_),
    .B2(_15149_),
    .ZN(_02779_));
 NOR2_X1 _25767_ (.A1(_02331_),
    .A2(_02779_),
    .ZN(_02780_));
 AOI222_X2 _25768_ (.A1(_02742_),
    .A2(_02754_),
    .B1(_02761_),
    .B2(_02769_),
    .C1(_02774_),
    .C2(_02780_),
    .ZN(_00116_));
 NAND2_X1 _25769_ (.A1(_02396_),
    .A2(_02436_),
    .ZN(_02781_));
 NAND2_X1 _25770_ (.A1(_02379_),
    .A2(_02425_),
    .ZN(_02782_));
 NOR2_X4 _25771_ (.A1(_02711_),
    .A2(_02402_),
    .ZN(_02783_));
 NOR2_X4 _25772_ (.A1(_02783_),
    .A2(_02369_),
    .ZN(_02784_));
 AOI21_X1 _25773_ (.A(_02707_),
    .B1(_02523_),
    .B2(_02317_),
    .ZN(_02785_));
 AOI221_X2 _25774_ (.A(_02325_),
    .B1(_02784_),
    .B2(_02782_),
    .C1(_02785_),
    .C2(_02383_),
    .ZN(_02786_));
 OR2_X1 _25775_ (.A1(_02379_),
    .A2(_02477_),
    .ZN(_02787_));
 NOR2_X2 _25776_ (.A1(_02453_),
    .A2(_02315_),
    .ZN(_02788_));
 AOI21_X1 _25777_ (.A(_02788_),
    .B1(_02318_),
    .B2(_02399_),
    .ZN(_02789_));
 OAI221_X1 _25778_ (.A(_02509_),
    .B1(_02690_),
    .B2(_02787_),
    .C1(_02789_),
    .C2(_02411_),
    .ZN(_02790_));
 OAI221_X1 _25779_ (.A(_02475_),
    .B1(_02344_),
    .B2(_02422_),
    .C1(_02404_),
    .C2(_02640_),
    .ZN(_02791_));
 OAI21_X1 _25780_ (.A(_02790_),
    .B1(_02791_),
    .B2(_02382_),
    .ZN(_02792_));
 AOI211_X2 _25781_ (.A(_02786_),
    .B(_02781_),
    .C1(_02792_),
    .C2(_02447_),
    .ZN(_02793_));
 AND2_X1 _25782_ (.A1(_02570_),
    .A2(_02667_),
    .ZN(_02794_));
 OAI221_X2 _25783_ (.A(_02509_),
    .B1(_02404_),
    .B2(_02374_),
    .C1(_02794_),
    .C2(_02313_),
    .ZN(_02795_));
 AOI221_X2 _25784_ (.A(_02361_),
    .B1(_02342_),
    .B2(_02629_),
    .C1(_02364_),
    .C2(_02453_),
    .ZN(_02796_));
 NOR2_X1 _25785_ (.A1(_02434_),
    .A2(_02796_),
    .ZN(_02797_));
 NOR2_X1 _25786_ (.A1(_02371_),
    .A2(_02315_),
    .ZN(_02798_));
 MUX2_X1 _25787_ (.A(_02788_),
    .B(_02798_),
    .S(_02349_),
    .Z(_02799_));
 NAND2_X1 _25788_ (.A1(_02390_),
    .A2(_02375_),
    .ZN(_02800_));
 AOI21_X1 _25789_ (.A(_02799_),
    .B1(_02542_),
    .B2(_02800_),
    .ZN(_02801_));
 INV_X1 _25790_ (.A(_02371_),
    .ZN(_02802_));
 OAI22_X2 _25791_ (.A1(_02802_),
    .A2(_02343_),
    .B1(_02579_),
    .B2(_02495_),
    .ZN(_02803_));
 MUX2_X1 _25792_ (.A(_02801_),
    .B(_02803_),
    .S(_02518_),
    .Z(_02804_));
 AOI221_X2 _25793_ (.A(_02587_),
    .B1(_02795_),
    .B2(_02797_),
    .C1(_02804_),
    .C2(_02435_),
    .ZN(_02805_));
 OAI221_X1 _25794_ (.A(_02603_),
    .B1(_02623_),
    .B2(_02385_),
    .C1(_02625_),
    .C2(_02707_),
    .ZN(_02806_));
 AND2_X1 _25795_ (.A1(_02403_),
    .A2(_02537_),
    .ZN(_02807_));
 AOI221_X1 _25796_ (.A(_02807_),
    .B1(_02484_),
    .B2(_02295_),
    .C1(_02483_),
    .C2(_02443_),
    .ZN(_02808_));
 OAI21_X1 _25797_ (.A(_02806_),
    .B1(_02808_),
    .B2(_02547_),
    .ZN(_02809_));
 AOI21_X1 _25798_ (.A(_15133_),
    .B1(_02344_),
    .B2(_02279_),
    .ZN(_02810_));
 OAI21_X1 _25799_ (.A(_02591_),
    .B1(_02669_),
    .B2(_02810_),
    .ZN(_02811_));
 OAI21_X1 _25800_ (.A(_02582_),
    .B1(_02579_),
    .B2(_02443_),
    .ZN(_02812_));
 OAI21_X1 _25801_ (.A(_02811_),
    .B1(_02812_),
    .B2(_02799_),
    .ZN(_02813_));
 NOR4_X2 _25802_ (.A1(_02414_),
    .A2(_02436_),
    .A3(_02809_),
    .A4(_02813_),
    .ZN(_02814_));
 NAND2_X1 _25803_ (.A1(_02414_),
    .A2(_02436_),
    .ZN(_02815_));
 NAND2_X1 _25804_ (.A1(_02362_),
    .A2(_02391_),
    .ZN(_02816_));
 NAND3_X1 _25805_ (.A1(_15133_),
    .A2(_02383_),
    .A3(_02344_),
    .ZN(_02817_));
 AOI21_X1 _25806_ (.A(net145),
    .B1(_02816_),
    .B2(_02817_),
    .ZN(_02818_));
 NOR3_X1 _25807_ (.A1(_02509_),
    .A2(_02411_),
    .A3(_02576_),
    .ZN(_02819_));
 AOI22_X1 _25808_ (.A1(net731),
    .A2(_02518_),
    .B1(_02376_),
    .B2(_02598_),
    .ZN(_02820_));
 OAI221_X1 _25809_ (.A(_02325_),
    .B1(_02458_),
    .B2(_02577_),
    .C1(_02820_),
    .C2(_15133_),
    .ZN(_02821_));
 NOR3_X1 _25810_ (.A1(_02818_),
    .A2(_02819_),
    .A3(_02821_),
    .ZN(_02822_));
 NAND2_X1 _25811_ (.A1(_02378_),
    .A2(_02411_),
    .ZN(_02823_));
 AOI21_X1 _25812_ (.A(_02636_),
    .B1(_02823_),
    .B2(_02678_),
    .ZN(_02824_));
 OAI21_X1 _25813_ (.A(_02582_),
    .B1(_02579_),
    .B2(net1044),
    .ZN(_02825_));
 NOR2_X1 _25814_ (.A1(_02824_),
    .A2(_02825_),
    .ZN(_02826_));
 MUX2_X1 _25815_ (.A(net1042),
    .B(_02407_),
    .S(_02349_),
    .Z(_02827_));
 AOI221_X2 _25816_ (.A(_02547_),
    .B1(_02827_),
    .B2(_02598_),
    .C1(_02483_),
    .C2(_02521_),
    .ZN(_02828_));
 NOR4_X1 _25817_ (.A1(_02815_),
    .A2(_02822_),
    .A3(_02826_),
    .A4(_02828_),
    .ZN(_02829_));
 OR4_X2 _25818_ (.A1(_02793_),
    .A2(_02805_),
    .A3(_02814_),
    .A4(_02829_),
    .ZN(_00117_));
 AOI221_X2 _25819_ (.A(_02370_),
    .B1(_02499_),
    .B2(_02699_),
    .C1(_02522_),
    .C2(_02636_),
    .ZN(_02830_));
 NOR2_X1 _25820_ (.A1(_02391_),
    .A2(_02719_),
    .ZN(_02831_));
 AOI221_X1 _25821_ (.A(_02363_),
    .B1(_02536_),
    .B2(_02831_),
    .C1(_02415_),
    .C2(_15144_),
    .ZN(_02832_));
 NOR2_X1 _25822_ (.A1(_02434_),
    .A2(_02436_),
    .ZN(_02833_));
 OAI221_X1 _25823_ (.A(_02449_),
    .B1(_02318_),
    .B2(_15122_),
    .C1(net580),
    .C2(_02579_),
    .ZN(_02834_));
 OAI221_X1 _25824_ (.A(_02439_),
    .B1(_02506_),
    .B2(_02344_),
    .C1(_02404_),
    .C2(_02374_),
    .ZN(_02835_));
 AOI21_X1 _25825_ (.A(net145),
    .B1(_02313_),
    .B2(_02762_),
    .ZN(_02836_));
 OAI221_X1 _25826_ (.A(_02833_),
    .B1(_02763_),
    .B2(_02834_),
    .C1(_02835_),
    .C2(_02836_),
    .ZN(_02837_));
 AOI21_X2 _25827_ (.A(net724),
    .B1(_02296_),
    .B2(_02279_),
    .ZN(_02838_));
 NOR2_X1 _25828_ (.A1(_15143_),
    .A2(_15152_),
    .ZN(_02839_));
 AOI221_X1 _25829_ (.A(_02621_),
    .B1(_02766_),
    .B2(_02838_),
    .C1(_02839_),
    .C2(_02375_),
    .ZN(_02840_));
 OR2_X1 _25830_ (.A1(_02331_),
    .A2(_02840_),
    .ZN(_02841_));
 OR2_X1 _25831_ (.A1(_15145_),
    .A2(_02375_),
    .ZN(_02842_));
 NAND2_X1 _25832_ (.A1(_02521_),
    .A2(_02317_),
    .ZN(_02843_));
 NAND3_X1 _25833_ (.A1(_02376_),
    .A2(_02614_),
    .A3(_02843_),
    .ZN(_02844_));
 NAND3_X1 _25834_ (.A1(_02356_),
    .A2(_02842_),
    .A3(_02844_),
    .ZN(_02845_));
 AOI21_X1 _25835_ (.A(_02548_),
    .B1(_02391_),
    .B2(_02378_),
    .ZN(_02846_));
 AOI211_X2 _25836_ (.A(_02402_),
    .B(_02729_),
    .C1(_02403_),
    .C2(_02407_),
    .ZN(_02847_));
 OAI21_X1 _25837_ (.A(_02395_),
    .B1(_02846_),
    .B2(_02847_),
    .ZN(_02848_));
 AND3_X1 _25838_ (.A1(_02475_),
    .A2(_02845_),
    .A3(_02848_),
    .ZN(_02849_));
 OR3_X2 _25839_ (.A1(_02471_),
    .A2(_02598_),
    .A3(_02646_),
    .ZN(_02850_));
 NAND2_X1 _25840_ (.A1(_02351_),
    .A2(_02567_),
    .ZN(_02851_));
 AOI21_X2 _25841_ (.A(_02363_),
    .B1(_02850_),
    .B2(_02851_),
    .ZN(_02852_));
 OAI33_X1 _25842_ (.A1(_02830_),
    .A2(_02832_),
    .A3(_02837_),
    .B1(_02852_),
    .B2(_02849_),
    .B3(_02841_),
    .ZN(_02853_));
 NOR2_X1 _25843_ (.A1(_02544_),
    .A2(_02644_),
    .ZN(_02854_));
 NOR2_X1 _25844_ (.A1(_02344_),
    .A2(_02666_),
    .ZN(_02855_));
 NOR3_X1 _25845_ (.A1(_02319_),
    .A2(_02392_),
    .A3(_02855_),
    .ZN(_02856_));
 OAI21_X1 _25846_ (.A(_02449_),
    .B1(_02854_),
    .B2(_02856_),
    .ZN(_02857_));
 AOI21_X1 _25847_ (.A(_02706_),
    .B1(_02416_),
    .B2(_15122_),
    .ZN(_02858_));
 OAI21_X1 _25848_ (.A(_02636_),
    .B1(_02415_),
    .B2(_02666_),
    .ZN(_02859_));
 NOR2_X1 _25849_ (.A1(_02552_),
    .A2(_02859_),
    .ZN(_02860_));
 OAI21_X1 _25850_ (.A(_02486_),
    .B1(_02858_),
    .B2(_02860_),
    .ZN(_02861_));
 AOI22_X1 _25851_ (.A1(_02495_),
    .A2(_02364_),
    .B1(_02483_),
    .B2(_02378_),
    .ZN(_02862_));
 AOI21_X2 _25852_ (.A(_02719_),
    .B1(_02316_),
    .B2(net1042),
    .ZN(_02863_));
 OR2_X1 _25853_ (.A1(_02400_),
    .A2(_02863_),
    .ZN(_02864_));
 NAND3_X1 _25854_ (.A1(_02439_),
    .A2(_02862_),
    .A3(_02864_),
    .ZN(_02865_));
 AOI21_X1 _25855_ (.A(_02646_),
    .B1(_02411_),
    .B2(_02802_),
    .ZN(_02866_));
 OAI221_X1 _25856_ (.A(_02510_),
    .B1(_02444_),
    .B2(net732),
    .C1(_02866_),
    .C2(_02319_),
    .ZN(_02867_));
 NAND4_X1 _25857_ (.A1(_02857_),
    .A2(_02861_),
    .A3(_02865_),
    .A4(_02867_),
    .ZN(_02868_));
 NAND2_X1 _25858_ (.A1(_02598_),
    .A2(_02762_),
    .ZN(_02869_));
 OAI21_X1 _25859_ (.A(_02506_),
    .B1(_02317_),
    .B2(net732),
    .ZN(_02870_));
 MUX2_X1 _25860_ (.A(_02539_),
    .B(_02870_),
    .S(_02343_),
    .Z(_02871_));
 AOI221_X1 _25861_ (.A(_02356_),
    .B1(_02784_),
    .B2(_02869_),
    .C1(_02871_),
    .C2(_02475_),
    .ZN(_02872_));
 MUX2_X1 _25862_ (.A(_02640_),
    .B(_02371_),
    .S(_02342_),
    .Z(_02873_));
 AOI221_X1 _25863_ (.A(_02362_),
    .B1(_02483_),
    .B2(net145),
    .C1(_02873_),
    .C2(_02598_),
    .ZN(_02874_));
 NOR3_X1 _25864_ (.A1(_02397_),
    .A2(_02595_),
    .A3(_02874_),
    .ZN(_02875_));
 OR2_X1 _25865_ (.A1(_02872_),
    .A2(_02875_),
    .ZN(_02876_));
 AOI221_X2 _25866_ (.A(_02853_),
    .B1(_02868_),
    .B2(_02438_),
    .C1(_02876_),
    .C2(_02448_),
    .ZN(_00118_));
 AOI21_X1 _25867_ (.A(_02426_),
    .B1(_02473_),
    .B2(_02678_),
    .ZN(_02877_));
 OR2_X1 _25868_ (.A1(_02558_),
    .A2(_02877_),
    .ZN(_02878_));
 OAI21_X1 _25869_ (.A(_02627_),
    .B1(_02317_),
    .B2(_02390_),
    .ZN(_02879_));
 MUX2_X1 _25870_ (.A(_15152_),
    .B(_02879_),
    .S(_02343_),
    .Z(_02880_));
 AOI21_X1 _25871_ (.A(_02447_),
    .B1(_02880_),
    .B2(_02509_),
    .ZN(_02881_));
 OAI221_X1 _25872_ (.A(_02509_),
    .B1(_02411_),
    .B2(_02443_),
    .C1(_02404_),
    .C2(_02332_),
    .ZN(_02882_));
 OR3_X1 _25873_ (.A1(_02636_),
    .A2(_02518_),
    .A3(_02583_),
    .ZN(_02883_));
 NAND4_X1 _25874_ (.A1(_02636_),
    .A2(_02475_),
    .A3(_02377_),
    .A4(_02513_),
    .ZN(_02884_));
 NAND3_X1 _25875_ (.A1(_02882_),
    .A2(_02883_),
    .A3(_02884_),
    .ZN(_02885_));
 AOI221_X1 _25876_ (.A(_02815_),
    .B1(_02878_),
    .B2(_02881_),
    .C1(_02885_),
    .C2(_02447_),
    .ZN(_02886_));
 NOR2_X1 _25877_ (.A1(_15129_),
    .A2(_02311_),
    .ZN(_02887_));
 OAI21_X1 _25878_ (.A(_02342_),
    .B1(_02425_),
    .B2(_02887_),
    .ZN(_02888_));
 OAI221_X2 _25879_ (.A(_02888_),
    .B1(_02526_),
    .B2(_02442_),
    .C1(_02405_),
    .C2(_02444_),
    .ZN(_02889_));
 OAI21_X1 _25880_ (.A(_02402_),
    .B1(_02403_),
    .B2(_02366_),
    .ZN(_02890_));
 OAI21_X2 _25881_ (.A(_02890_),
    .B1(_02755_),
    .B2(_02312_),
    .ZN(_02891_));
 AOI221_X2 _25882_ (.A(_02330_),
    .B1(_02603_),
    .B2(_02889_),
    .C1(_02891_),
    .C2(_02591_),
    .ZN(_02892_));
 NOR2_X1 _25883_ (.A1(_02369_),
    .A2(_02349_),
    .ZN(_02893_));
 AND3_X1 _25884_ (.A1(_02361_),
    .A2(_02349_),
    .A3(_02506_),
    .ZN(_02894_));
 AOI221_X2 _25885_ (.A(_02324_),
    .B1(_02893_),
    .B2(_02863_),
    .C1(_02894_),
    .C2(_02476_),
    .ZN(_02895_));
 AOI222_X2 _25886_ (.A1(_15122_),
    .A2(_02430_),
    .B1(_02483_),
    .B2(_02453_),
    .C1(_02521_),
    .C2(_02484_),
    .ZN(_02896_));
 OAI21_X1 _25887_ (.A(_02895_),
    .B1(_02896_),
    .B2(_02509_),
    .ZN(_02897_));
 NAND3_X1 _25888_ (.A1(_02312_),
    .A2(_02639_),
    .A3(_02643_),
    .ZN(_02898_));
 AOI21_X1 _25889_ (.A(_02898_),
    .B1(_02376_),
    .B2(_02495_),
    .ZN(_02899_));
 AOI21_X1 _25890_ (.A(_02598_),
    .B1(_02380_),
    .B2(_02609_),
    .ZN(_02900_));
 AOI21_X1 _25891_ (.A(_02899_),
    .B1(_02900_),
    .B2(_02473_),
    .ZN(_02901_));
 OAI21_X1 _25892_ (.A(_02318_),
    .B1(_02380_),
    .B2(_02407_),
    .ZN(_02902_));
 OAI22_X1 _25893_ (.A1(_02624_),
    .A2(_02902_),
    .B1(_02705_),
    .B2(_02636_),
    .ZN(_02903_));
 AOI22_X2 _25894_ (.A1(_02603_),
    .A2(_02901_),
    .B1(_02903_),
    .B2(_02591_),
    .ZN(_02904_));
 NAND2_X1 _25895_ (.A1(_02766_),
    .A2(_02838_),
    .ZN(_02905_));
 NOR2_X1 _25896_ (.A1(_02605_),
    .A2(_02535_),
    .ZN(_02906_));
 OAI21_X1 _25897_ (.A(_02402_),
    .B1(_02350_),
    .B2(_02378_),
    .ZN(_02907_));
 OAI22_X1 _25898_ (.A1(_02405_),
    .A2(_02312_),
    .B1(_02563_),
    .B2(_02907_),
    .ZN(_02908_));
 INV_X1 _25899_ (.A(_02547_),
    .ZN(_02909_));
 AOI221_X2 _25900_ (.A(_02504_),
    .B1(_02905_),
    .B2(_02906_),
    .C1(_02908_),
    .C2(_02909_),
    .ZN(_02910_));
 AOI221_X2 _25901_ (.A(_02414_),
    .B1(_02892_),
    .B2(_02897_),
    .C1(_02904_),
    .C2(_02910_),
    .ZN(_02911_));
 OAI21_X2 _25902_ (.A(_02318_),
    .B1(_02471_),
    .B2(_02707_),
    .ZN(_02912_));
 AOI21_X1 _25903_ (.A(_02518_),
    .B1(_02430_),
    .B2(_02443_),
    .ZN(_02913_));
 AOI21_X1 _25904_ (.A(_02684_),
    .B1(_02400_),
    .B2(_02443_),
    .ZN(_02914_));
 AOI221_X2 _25905_ (.A(_02447_),
    .B1(_02912_),
    .B2(_02913_),
    .C1(_02914_),
    .C2(_02800_),
    .ZN(_02915_));
 NAND4_X1 _25906_ (.A1(_02495_),
    .A2(_02598_),
    .A3(_02362_),
    .A4(_02343_),
    .ZN(_02916_));
 NAND4_X1 _25907_ (.A1(_15122_),
    .A2(_02548_),
    .A3(_02383_),
    .A4(_02391_),
    .ZN(_02917_));
 NAND3_X1 _25908_ (.A1(_02325_),
    .A2(_02916_),
    .A3(_02917_),
    .ZN(_02918_));
 NAND2_X1 _25909_ (.A1(_02383_),
    .A2(_02343_),
    .ZN(_02919_));
 OAI21_X1 _25910_ (.A(_02919_),
    .B1(_02816_),
    .B2(net1044),
    .ZN(_02920_));
 OAI21_X1 _25911_ (.A(_02526_),
    .B1(_02577_),
    .B2(_02313_),
    .ZN(_02921_));
 AOI221_X2 _25912_ (.A(_02918_),
    .B1(_02920_),
    .B2(_15133_),
    .C1(_02921_),
    .C2(net1044),
    .ZN(_02922_));
 NOR3_X1 _25913_ (.A1(_02915_),
    .A2(_02587_),
    .A3(_02922_),
    .ZN(_02923_));
 OR3_X2 _25914_ (.A1(_02923_),
    .A2(_02911_),
    .A3(_02886_),
    .ZN(_00119_));
 INV_X1 _25915_ (.A(\u0.tmp_w[9] ),
    .ZN(_02924_));
 NOR2_X1 _25916_ (.A1(_02924_),
    .A2(_09823_),
    .ZN(_02925_));
 NOR2_X1 _25917_ (.A1(\u0.tmp_w[9] ),
    .A2(_09823_),
    .ZN(_02926_));
 XNOR2_X2 _25918_ (.A(net974),
    .B(net658),
    .ZN(_02927_));
 XNOR2_X2 _25919_ (.A(_02927_),
    .B(_11185_),
    .ZN(_02928_));
 XNOR2_X1 _25920_ (.A(_11136_),
    .B(_11135_),
    .ZN(_02929_));
 XNOR2_X1 _25921_ (.A(_11114_),
    .B(_02929_),
    .ZN(_02930_));
 XNOR2_X2 _25922_ (.A(_02930_),
    .B(_02928_),
    .ZN(_02931_));
 MUX2_X1 _25923_ (.A(_02925_),
    .B(_02926_),
    .S(_02931_),
    .Z(_02932_));
 NAND3_X1 _25924_ (.A1(net1049),
    .A2(_09135_),
    .A3(_00473_),
    .ZN(_02933_));
 NAND2_X1 _25925_ (.A1(_02924_),
    .A2(_09135_),
    .ZN(_02934_));
 OAI21_X2 _25926_ (.A(_02933_),
    .B1(_02934_),
    .B2(_00473_),
    .ZN(_02935_));
 NOR2_X4 _25927_ (.A1(_02932_),
    .A2(_02935_),
    .ZN(_02936_));
 INV_X8 _25928_ (.A(net884),
    .ZN(_02937_));
 OAI21_X4 clone270 (.A(net10),
    .B1(_11231_),
    .B2(_11235_),
    .ZN(net733));
 BUF_X16 _25930_ (.A(_02937_),
    .Z(_15164_));
 XNOR2_X1 _25931_ (.A(_11135_),
    .B(_11117_),
    .ZN(_02939_));
 XOR2_X1 _25932_ (.A(_11183_),
    .B(_11184_),
    .Z(_02940_));
 NAND3_X4 _25933_ (.A1(_11191_),
    .A2(_06457_),
    .A3(_02940_),
    .ZN(_02941_));
 NOR2_X1 _25934_ (.A1(_06457_),
    .A2(_11938_),
    .ZN(_02942_));
 NAND2_X1 _25935_ (.A1(_11185_),
    .A2(_02942_),
    .ZN(_02943_));
 AOI21_X4 _25936_ (.A(_02939_),
    .B1(_02941_),
    .B2(_02943_),
    .ZN(_02944_));
 XOR2_X1 _25937_ (.A(_11135_),
    .B(_11117_),
    .Z(_02945_));
 NAND2_X1 _25938_ (.A1(_02940_),
    .A2(_02942_),
    .ZN(_02946_));
 NAND3_X1 _25939_ (.A1(_06457_),
    .A2(_09116_),
    .A3(_11185_),
    .ZN(_02947_));
 AOI21_X1 _25940_ (.A(_02945_),
    .B1(_02946_),
    .B2(_02947_),
    .ZN(_02948_));
 INV_X1 _25941_ (.A(_06457_),
    .ZN(_02949_));
 NAND3_X1 _25942_ (.A1(_02949_),
    .A2(_09103_),
    .A3(_00474_),
    .ZN(_02950_));
 NAND2_X1 _25943_ (.A1(_06457_),
    .A2(_09103_),
    .ZN(_02951_));
 OAI21_X1 _25944_ (.A(_02950_),
    .B1(_02951_),
    .B2(_00474_),
    .ZN(_02952_));
 OR3_X4 _25945_ (.A1(_02948_),
    .A2(_02944_),
    .A3(_02952_),
    .ZN(_02953_));
 BUF_X16 _25946_ (.A(_02953_),
    .Z(_02954_));
 INV_X8 _25947_ (.A(_02954_),
    .ZN(_02955_));
 BUF_X8 _25948_ (.A(_02955_),
    .Z(_15169_));
 XNOR2_X1 _25949_ (.A(_11158_),
    .B(_13864_),
    .ZN(_02956_));
 OR3_X1 _25950_ (.A1(_06491_),
    .A2(_09030_),
    .A3(net959),
    .ZN(_02957_));
 NAND3_X1 _25951_ (.A1(_06491_),
    .A2(_09195_),
    .A3(net959),
    .ZN(_02958_));
 AOI21_X2 _25952_ (.A(_02956_),
    .B1(_02957_),
    .B2(_02958_),
    .ZN(_02959_));
 XNOR2_X1 _25953_ (.A(_11158_),
    .B(_13862_),
    .ZN(_02960_));
 OR3_X1 _25954_ (.A1(_06479_),
    .A2(_09727_),
    .A3(net959),
    .ZN(_02961_));
 NAND3_X1 _25955_ (.A1(_06479_),
    .A2(net1085),
    .A3(net959),
    .ZN(_02962_));
 AOI21_X2 _25956_ (.A(_02960_),
    .B1(_02961_),
    .B2(_02962_),
    .ZN(_02963_));
 NAND3_X1 _25957_ (.A1(_06491_),
    .A2(_09730_),
    .A3(_00475_),
    .ZN(_02964_));
 NAND2_X1 _25958_ (.A1(_06479_),
    .A2(_09730_),
    .ZN(_02965_));
 OAI21_X2 _25959_ (.A(_02964_),
    .B1(_02965_),
    .B2(_00475_),
    .ZN(_02966_));
 NOR3_X4 _25960_ (.A1(_02966_),
    .A2(_02963_),
    .A3(_02959_),
    .ZN(_02967_));
 INV_X4 _25961_ (.A(net1037),
    .ZN(_02968_));
 BUF_X4 _25962_ (.A(_02968_),
    .Z(_02969_));
 BUF_X4 _25963_ (.A(_02969_),
    .Z(_02970_));
 BUF_X4 _25964_ (.A(_02970_),
    .Z(_02971_));
 BUF_X4 _25965_ (.A(_02971_),
    .Z(_15185_));
 BUF_X8 _25966_ (.A(_02936_),
    .Z(_02972_));
 BUF_X16 _25967_ (.A(_02972_),
    .Z(_15159_));
 BUF_X4 _25968_ (.A(net1037),
    .Z(_02973_));
 BUF_X4 _25969_ (.A(_02973_),
    .Z(_02974_));
 BUF_X4 _25970_ (.A(_02974_),
    .Z(_02975_));
 BUF_X4 _25971_ (.A(_02975_),
    .Z(_15178_));
 BUF_X8 _25972_ (.A(_15176_),
    .Z(_02976_));
 NAND2_X1 _25973_ (.A1(_11841_),
    .A2(\text_in_r[11] ),
    .ZN(_02977_));
 NAND3_X2 _25974_ (.A1(_06517_),
    .A2(_08975_),
    .A3(_02977_),
    .ZN(_02978_));
 OR2_X1 _25975_ (.A1(_06517_),
    .A2(_02977_),
    .ZN(_02979_));
 AND2_X1 _25976_ (.A1(_02978_),
    .A2(_02979_),
    .ZN(_02980_));
 BUF_X4 _25977_ (.A(_02980_),
    .Z(_02981_));
 BUF_X8 _25978_ (.A(_02981_),
    .Z(_02982_));
 NAND2_X1 _25979_ (.A1(_06517_),
    .A2(_02977_),
    .ZN(_02983_));
 OR2_X1 _25980_ (.A1(_06517_),
    .A2(_00991_),
    .ZN(_02984_));
 XNOR2_X1 _25981_ (.A(_11245_),
    .B(_11184_),
    .ZN(_02985_));
 XNOR2_X1 _25982_ (.A(_11164_),
    .B(_11223_),
    .ZN(_02986_));
 XNOR2_X2 _25983_ (.A(_02985_),
    .B(_02986_),
    .ZN(_02987_));
 XNOR2_X1 _25984_ (.A(_11183_),
    .B(_13930_),
    .ZN(_02988_));
 XNOR2_X2 _25985_ (.A(_02987_),
    .B(_02988_),
    .ZN(_02989_));
 MUX2_X2 _25986_ (.A(_02983_),
    .B(_02984_),
    .S(_02989_),
    .Z(_02990_));
 BUF_X8 _25987_ (.A(_02990_),
    .Z(_02991_));
 AOI21_X4 _25988_ (.A(_02976_),
    .B1(_02982_),
    .B2(_02991_),
    .ZN(_02992_));
 NAND2_X4 _25989_ (.A1(_02978_),
    .A2(_02979_),
    .ZN(_02993_));
 AND2_X1 _25990_ (.A1(_06517_),
    .A2(_02977_),
    .ZN(_02994_));
 NOR2_X1 _25991_ (.A1(_06517_),
    .A2(_08975_),
    .ZN(_02995_));
 MUX2_X2 _25992_ (.A(_02994_),
    .B(_02995_),
    .S(_02989_),
    .Z(_02996_));
 NOR2_X4 _25993_ (.A1(_02993_),
    .A2(_02996_),
    .ZN(_02997_));
 BUF_X4 _25994_ (.A(_02997_),
    .Z(_02998_));
 BUF_X4 _25995_ (.A(_02998_),
    .Z(_02999_));
 BUF_X4 _25996_ (.A(net884),
    .Z(_03000_));
 AOI211_X2 _25997_ (.A(_02970_),
    .B(_02992_),
    .C1(_02999_),
    .C2(_03000_),
    .ZN(_03001_));
 BUF_X8 clone200 (.A(_12606_),
    .Z(net200));
 BUF_X8 _25999_ (.A(_02993_),
    .Z(_03003_));
 BUF_X8 _26000_ (.A(_02996_),
    .Z(_03004_));
 NOR3_X4 _26001_ (.A1(net514),
    .A2(_03003_),
    .A3(_03004_),
    .ZN(_03005_));
 AOI21_X2 _26002_ (.A(_02954_),
    .B1(_02982_),
    .B2(_02991_),
    .ZN(_03006_));
 OR2_X1 _26003_ (.A1(_03005_),
    .A2(_03006_),
    .ZN(_03007_));
 AOI21_X1 _26004_ (.A(_03001_),
    .B1(_03007_),
    .B2(_15185_),
    .ZN(_03008_));
 XNOR2_X1 _26005_ (.A(_11265_),
    .B(_11184_),
    .ZN(_03009_));
 XNOR2_X1 _26006_ (.A(_11225_),
    .B(_11249_),
    .ZN(_03010_));
 XNOR2_X2 _26007_ (.A(_03009_),
    .B(_03010_),
    .ZN(_03011_));
 XNOR2_X1 _26008_ (.A(_13914_),
    .B(_03011_),
    .ZN(_03012_));
 MUX2_X2 _26009_ (.A(\text_in_r[12] ),
    .B(_03012_),
    .S(_09075_),
    .Z(_03013_));
 XNOR2_X2 _26010_ (.A(_06533_),
    .B(_03013_),
    .ZN(_03014_));
 BUF_X4 _26011_ (.A(_03014_),
    .Z(_03015_));
 XOR2_X2 _26012_ (.A(_11246_),
    .B(_11262_),
    .Z(_03016_));
 NAND3_X1 _26013_ (.A1(_06546_),
    .A2(_09175_),
    .A3(_03016_),
    .ZN(_03017_));
 NOR2_X1 _26014_ (.A1(_06546_),
    .A2(_09179_),
    .ZN(_03018_));
 NAND2_X1 _26015_ (.A1(_03016_),
    .A2(_03018_),
    .ZN(_03019_));
 XNOR2_X2 _26016_ (.A(_11250_),
    .B(_11203_),
    .ZN(_03020_));
 MUX2_X1 _26017_ (.A(_03017_),
    .B(_03019_),
    .S(_03020_),
    .Z(_03021_));
 XNOR2_X1 _26018_ (.A(_11246_),
    .B(_11262_),
    .ZN(_03022_));
 NAND2_X1 _26019_ (.A1(_03022_),
    .A2(_03018_),
    .ZN(_03023_));
 NAND3_X1 _26020_ (.A1(_06546_),
    .A2(_09076_),
    .A3(_03022_),
    .ZN(_03024_));
 MUX2_X1 _26021_ (.A(_03023_),
    .B(_03024_),
    .S(_03020_),
    .Z(_03025_));
 OR3_X2 _26022_ (.A1(_06546_),
    .A2(_09138_),
    .A3(\text_in_r[13] ),
    .ZN(_03026_));
 NAND3_X2 _26023_ (.A1(_06546_),
    .A2(_09824_),
    .A3(\text_in_r[13] ),
    .ZN(_03027_));
 AND4_X1 _26024_ (.A1(_03021_),
    .A2(_03025_),
    .A3(_03026_),
    .A4(_03027_),
    .ZN(_03028_));
 BUF_X4 _26025_ (.A(_03028_),
    .Z(_03029_));
 NOR2_X4 _26026_ (.A1(_03015_),
    .A2(_03029_),
    .ZN(_03030_));
 NAND4_X4 _26027_ (.A1(_03021_),
    .A2(_03025_),
    .A3(_03026_),
    .A4(_03027_),
    .ZN(_03031_));
 BUF_X4 _26028_ (.A(_03031_),
    .Z(_03032_));
 NOR2_X2 _26029_ (.A1(_03015_),
    .A2(_03032_),
    .ZN(_03033_));
 CLKBUF_X3 _26030_ (.A(_02975_),
    .Z(_03034_));
 NOR3_X4 _26031_ (.A1(_02955_),
    .A2(_03003_),
    .A3(_03004_),
    .ZN(_03035_));
 BUF_X4 _26032_ (.A(_15161_),
    .Z(_03036_));
 AOI21_X4 _26033_ (.A(_03036_),
    .B1(_02982_),
    .B2(_02991_),
    .ZN(_03037_));
 OAI21_X1 _26034_ (.A(_03034_),
    .B1(_03035_),
    .B2(_03037_),
    .ZN(_03038_));
 BUF_X4 _26035_ (.A(_02997_),
    .Z(_03039_));
 AOI21_X1 _26036_ (.A(_02992_),
    .B1(_03039_),
    .B2(net515),
    .ZN(_03040_));
 OAI21_X1 _26037_ (.A(_03038_),
    .B1(_03040_),
    .B2(_15178_),
    .ZN(_03041_));
 AOI22_X1 _26038_ (.A1(_03008_),
    .A2(_03030_),
    .B1(_03033_),
    .B2(_03041_),
    .ZN(_03042_));
 XOR2_X2 _26039_ (.A(_06533_),
    .B(_03013_),
    .Z(_03043_));
 BUF_X4 _26040_ (.A(_03043_),
    .Z(_03044_));
 NOR2_X4 _26041_ (.A1(_03044_),
    .A2(_03032_),
    .ZN(_03045_));
 BUF_X4 _26042_ (.A(_02982_),
    .Z(_03046_));
 BUF_X4 _26043_ (.A(_02991_),
    .Z(_03047_));
 NAND3_X4 _26044_ (.A1(net1084),
    .A2(_03046_),
    .A3(_03047_),
    .ZN(_03048_));
 BUF_X4 _26045_ (.A(_03003_),
    .Z(_03049_));
 BUF_X4 _26046_ (.A(_03004_),
    .Z(_03050_));
 OAI21_X2 _26047_ (.A(net515),
    .B1(_03049_),
    .B2(_03050_),
    .ZN(_03051_));
 AOI21_X1 _26048_ (.A(_15178_),
    .B1(_03048_),
    .B2(_03051_),
    .ZN(_03052_));
 BUF_X8 _26049_ (.A(_15167_),
    .Z(_03053_));
 OAI21_X4 _26050_ (.A(_02973_),
    .B1(_03003_),
    .B2(_03004_),
    .ZN(_03054_));
 NOR2_X1 _26051_ (.A1(_03053_),
    .A2(_03054_),
    .ZN(_03055_));
 OAI21_X1 _26052_ (.A(_03045_),
    .B1(_03052_),
    .B2(_03055_),
    .ZN(_03056_));
 XNOR2_X1 _26053_ (.A(_11263_),
    .B(_13904_),
    .ZN(_03057_));
 XNOR2_X1 _26054_ (.A(_11186_),
    .B(_03057_),
    .ZN(_03058_));
 MUX2_X2 _26055_ (.A(\text_in_r[14] ),
    .B(_03058_),
    .S(_09803_),
    .Z(_03059_));
 XOR2_X2 _26056_ (.A(_06554_),
    .B(_03059_),
    .Z(_03060_));
 XNOR2_X1 _26057_ (.A(_11198_),
    .B(_11184_),
    .ZN(_03061_));
 XNOR2_X1 _26058_ (.A(_11121_),
    .B(_03061_),
    .ZN(_03062_));
 XNOR2_X1 _26059_ (.A(_11199_),
    .B(_03062_),
    .ZN(_03063_));
 MUX2_X2 _26060_ (.A(\text_in_r[15] ),
    .B(_03063_),
    .S(_10571_),
    .Z(_03064_));
 XNOR2_X2 _26061_ (.A(_06563_),
    .B(_03064_),
    .ZN(_03065_));
 NAND2_X2 _26062_ (.A1(_03060_),
    .A2(_03065_),
    .ZN(_03066_));
 INV_X1 _26063_ (.A(_03066_),
    .ZN(_03067_));
 NAND2_X1 _26064_ (.A1(_02981_),
    .A2(_02990_),
    .ZN(_03068_));
 BUF_X4 _26065_ (.A(_03068_),
    .Z(_03069_));
 BUF_X4 _26066_ (.A(_03069_),
    .Z(_03070_));
 BUF_X4 _26067_ (.A(_15174_),
    .Z(_03071_));
 INV_X2 _26068_ (.A(_03071_),
    .ZN(_03072_));
 MUX2_X1 _26069_ (.A(_03072_),
    .B(_02955_),
    .S(_02968_),
    .Z(_03073_));
 AOI21_X2 _26070_ (.A(_03044_),
    .B1(_03070_),
    .B2(_03073_),
    .ZN(_03074_));
 INV_X1 _26071_ (.A(_03074_),
    .ZN(_03075_));
 BUF_X4 _26072_ (.A(_03032_),
    .Z(_03076_));
 CLKBUF_X3 _26073_ (.A(_03076_),
    .Z(_03077_));
 NOR2_X2 _26074_ (.A1(_15159_),
    .A2(_02975_),
    .ZN(_03078_));
 CLKBUF_X3 _26075_ (.A(_03039_),
    .Z(_03079_));
 BUF_X8 _26076_ (.A(_15162_),
    .Z(_03080_));
 OAI21_X1 _26077_ (.A(_03079_),
    .B1(_02971_),
    .B2(net1045),
    .ZN(_03081_));
 OAI21_X1 _26078_ (.A(_03077_),
    .B1(_03078_),
    .B2(_03081_),
    .ZN(_03082_));
 OR2_X1 _26079_ (.A1(_03075_),
    .A2(_03082_),
    .ZN(_03083_));
 NAND4_X2 _26080_ (.A1(_03042_),
    .A2(_03056_),
    .A3(_03067_),
    .A4(_03083_),
    .ZN(_03084_));
 NOR2_X4 _26081_ (.A1(_03060_),
    .A2(_03065_),
    .ZN(_03085_));
 BUF_X4 _26082_ (.A(_03029_),
    .Z(_03086_));
 BUF_X4 _26083_ (.A(_03086_),
    .Z(_03087_));
 CLKBUF_X3 _26084_ (.A(_03087_),
    .Z(_03088_));
 BUF_X4 _26085_ (.A(_03044_),
    .Z(_03089_));
 BUF_X4 _26086_ (.A(_03089_),
    .Z(_03090_));
 AOI21_X1 _26087_ (.A(_03005_),
    .B1(_03070_),
    .B2(net1045),
    .ZN(_03091_));
 BUF_X4 _26088_ (.A(_02970_),
    .Z(_03092_));
 NAND3_X4 _26089_ (.A1(_02968_),
    .A2(_02981_),
    .A3(_02990_),
    .ZN(_03093_));
 BUF_X4 _26090_ (.A(_15170_),
    .Z(_03094_));
 OAI221_X1 _26091_ (.A(_03090_),
    .B1(_03091_),
    .B2(_03092_),
    .C1(_03093_),
    .C2(_03094_),
    .ZN(_03095_));
 CLKBUF_X3 _26092_ (.A(_03015_),
    .Z(_03096_));
 CLKBUF_X3 _26093_ (.A(_03096_),
    .Z(_03097_));
 INV_X4 _26094_ (.A(_15165_),
    .ZN(_03098_));
 AOI21_X4 _26095_ (.A(_03098_),
    .B1(_02981_),
    .B2(_02990_),
    .ZN(_03099_));
 NOR3_X4 _26096_ (.A1(_15162_),
    .A2(_02993_),
    .A3(_02996_),
    .ZN(_03100_));
 OR2_X1 _26097_ (.A1(_03099_),
    .A2(_03100_),
    .ZN(_03101_));
 OAI21_X4 _26098_ (.A(_02968_),
    .B1(_03003_),
    .B2(_03004_),
    .ZN(_03102_));
 BUF_X2 clone202 (.A(net203),
    .Z(net202));
 INV_X2 _26100_ (.A(net564),
    .ZN(_03104_));
 OAI221_X1 _26101_ (.A(_03097_),
    .B1(_03101_),
    .B2(_03092_),
    .C1(_03102_),
    .C2(_03104_),
    .ZN(_03105_));
 AND3_X1 _26102_ (.A1(_03088_),
    .A2(_03095_),
    .A3(_03105_),
    .ZN(_03106_));
 BUF_X4 _26103_ (.A(_03086_),
    .Z(_03107_));
 BUF_X4 _26104_ (.A(_15160_),
    .Z(_03108_));
 AOI21_X2 _26105_ (.A(_03108_),
    .B1(_02982_),
    .B2(_02991_),
    .ZN(_03109_));
 OAI21_X1 _26106_ (.A(_02974_),
    .B1(_03005_),
    .B2(_03109_),
    .ZN(_03110_));
 NOR3_X4 _26107_ (.A1(net1038),
    .A2(_03003_),
    .A3(_03004_),
    .ZN(_03111_));
 AOI21_X1 _26108_ (.A(_03044_),
    .B1(_03111_),
    .B2(_03053_),
    .ZN(_03112_));
 AND2_X1 _26109_ (.A1(_03110_),
    .A2(_03112_),
    .ZN(_03113_));
 BUF_X4 _26110_ (.A(_02969_),
    .Z(_03114_));
 BUF_X4 _26111_ (.A(_03114_),
    .Z(_03115_));
 OAI21_X4 _26112_ (.A(_02955_),
    .B1(_03003_),
    .B2(_03004_),
    .ZN(_03116_));
 CLKBUF_X3 _26113_ (.A(_03069_),
    .Z(_03117_));
 INV_X2 _26114_ (.A(_03080_),
    .ZN(_03118_));
 OAI21_X1 _26115_ (.A(_03116_),
    .B1(_03117_),
    .B2(_03118_),
    .ZN(_03119_));
 NAND2_X1 _26116_ (.A1(_03115_),
    .A2(_03119_),
    .ZN(_03120_));
 BUF_X4 _26117_ (.A(_03070_),
    .Z(_03121_));
 BUF_X8 _26118_ (.A(_03036_),
    .Z(_03122_));
 AOI22_X1 _26119_ (.A1(_15183_),
    .A2(_03121_),
    .B1(_03111_),
    .B2(_03122_),
    .ZN(_03123_));
 AOI221_X1 _26120_ (.A(_03107_),
    .B1(_03113_),
    .B2(_03120_),
    .C1(_03123_),
    .C2(_03090_),
    .ZN(_03124_));
 OAI21_X1 _26121_ (.A(_03085_),
    .B1(_03106_),
    .B2(_03124_),
    .ZN(_03125_));
 NAND2_X2 _26122_ (.A1(_02972_),
    .A2(net1084),
    .ZN(_03126_));
 NAND2_X2 _26123_ (.A1(_02955_),
    .A2(_02973_),
    .ZN(_03127_));
 AOI221_X2 _26124_ (.A(_03032_),
    .B1(_03126_),
    .B2(_03127_),
    .C1(_03039_),
    .C2(_03089_),
    .ZN(_03128_));
 NOR2_X1 _26125_ (.A1(_03015_),
    .A2(_02997_),
    .ZN(_03129_));
 NOR2_X2 _26126_ (.A1(net725),
    .A2(_02974_),
    .ZN(_03130_));
 INV_X1 _26127_ (.A(_03130_),
    .ZN(_03131_));
 OAI21_X1 _26128_ (.A(_03129_),
    .B1(_03131_),
    .B2(_03107_),
    .ZN(_03132_));
 INV_X4 _26129_ (.A(_03036_),
    .ZN(_03133_));
 BUF_X4 _26130_ (.A(_02969_),
    .Z(_03134_));
 NOR3_X1 _26131_ (.A1(_03133_),
    .A2(_03134_),
    .A3(_03086_),
    .ZN(_03135_));
 NOR3_X1 _26132_ (.A1(_03096_),
    .A2(_03121_),
    .A3(_03135_),
    .ZN(_03136_));
 BUF_X16 _26133_ (.A(_02954_),
    .Z(_15158_));
 AOI21_X1 _26134_ (.A(_03115_),
    .B1(_03087_),
    .B2(_15158_),
    .ZN(_03137_));
 NAND2_X1 _26135_ (.A1(_15169_),
    .A2(_03029_),
    .ZN(_03138_));
 OAI221_X1 _26136_ (.A(_03136_),
    .B1(_03137_),
    .B2(_15159_),
    .C1(_03034_),
    .C2(_03138_),
    .ZN(_03139_));
 AOI21_X1 _26137_ (.A(_03128_),
    .B1(_03132_),
    .B2(_03139_),
    .ZN(_03140_));
 XNOR2_X2 _26138_ (.A(_06554_),
    .B(_03059_),
    .ZN(_03141_));
 NAND2_X2 _26139_ (.A1(_03141_),
    .A2(_03065_),
    .ZN(_03142_));
 BUF_X4 _26140_ (.A(_03134_),
    .Z(_03143_));
 AOI21_X4 _26141_ (.A(_03094_),
    .B1(_02981_),
    .B2(_02990_),
    .ZN(_03144_));
 NOR3_X4 _26142_ (.A1(_03133_),
    .A2(_03049_),
    .A3(_03050_),
    .ZN(_03145_));
 NOR3_X1 _26143_ (.A1(_03143_),
    .A2(_03144_),
    .A3(_03145_),
    .ZN(_03146_));
 NOR3_X4 _26144_ (.A1(_03071_),
    .A2(_03003_),
    .A3(_03004_),
    .ZN(_03147_));
 NOR3_X1 _26145_ (.A1(_02975_),
    .A2(_03109_),
    .A3(_03147_),
    .ZN(_03148_));
 OAI21_X1 _26146_ (.A(_03045_),
    .B1(_03146_),
    .B2(_03148_),
    .ZN(_03149_));
 NOR2_X1 _26147_ (.A1(_03122_),
    .A2(_03054_),
    .ZN(_03150_));
 NAND3_X4 _26148_ (.A1(_02973_),
    .A2(_02982_),
    .A3(_02991_),
    .ZN(_03151_));
 NAND2_X1 _26149_ (.A1(_03102_),
    .A2(_03151_),
    .ZN(_03152_));
 AOI221_X1 _26150_ (.A(_03150_),
    .B1(_03152_),
    .B2(_03108_),
    .C1(_03094_),
    .C2(_03111_),
    .ZN(_03153_));
 NAND2_X4 _26151_ (.A1(_03014_),
    .A2(_03031_),
    .ZN(_03154_));
 OAI21_X1 _26152_ (.A(_03149_),
    .B1(_03154_),
    .B2(_03153_),
    .ZN(_03155_));
 OR3_X2 _26153_ (.A1(_03155_),
    .A2(_03142_),
    .A3(_03140_),
    .ZN(_03156_));
 BUF_X4 _26154_ (.A(_02973_),
    .Z(_03157_));
 AOI21_X4 _26155_ (.A(_03053_),
    .B1(_02982_),
    .B2(_02991_),
    .ZN(_03158_));
 OAI21_X2 _26156_ (.A(_03157_),
    .B1(_03100_),
    .B2(_03158_),
    .ZN(_03159_));
 AOI21_X1 _26157_ (.A(_03015_),
    .B1(_03111_),
    .B2(_03108_),
    .ZN(_03160_));
 OAI21_X1 _26158_ (.A(_03116_),
    .B1(_03069_),
    .B2(_02937_),
    .ZN(_03161_));
 NOR3_X2 _26159_ (.A1(_03036_),
    .A2(_03003_),
    .A3(_03004_),
    .ZN(_03162_));
 OR2_X1 _26160_ (.A1(_03144_),
    .A2(_03162_),
    .ZN(_03163_));
 MUX2_X1 _26161_ (.A(_03161_),
    .B(_03163_),
    .S(_03114_),
    .Z(_03164_));
 AOI221_X2 _26162_ (.A(_03076_),
    .B1(_03159_),
    .B2(_03160_),
    .C1(_03164_),
    .C2(_03096_),
    .ZN(_03165_));
 XOR2_X2 _26163_ (.A(_06563_),
    .B(_03064_),
    .Z(_03166_));
 NAND2_X1 _26164_ (.A1(_03060_),
    .A2(_03166_),
    .ZN(_03167_));
 AOI21_X4 _26165_ (.A(_02955_),
    .B1(_03046_),
    .B2(_03047_),
    .ZN(_03168_));
 NAND2_X1 _26166_ (.A1(_03015_),
    .A2(_03168_),
    .ZN(_03169_));
 NOR3_X4 _26167_ (.A1(net537),
    .A2(_02993_),
    .A3(_02996_),
    .ZN(_03170_));
 NOR2_X1 _26168_ (.A1(_03157_),
    .A2(_03170_),
    .ZN(_03171_));
 OAI21_X4 _26169_ (.A(net725),
    .B1(_03049_),
    .B2(_03050_),
    .ZN(_03172_));
 NAND3_X2 _26170_ (.A1(_15172_),
    .A2(_02982_),
    .A3(_02991_),
    .ZN(_03173_));
 AOI21_X1 _26171_ (.A(_02969_),
    .B1(_03172_),
    .B2(_03173_),
    .ZN(_03174_));
 OR2_X1 _26172_ (.A1(_03015_),
    .A2(_03174_),
    .ZN(_03175_));
 AOI221_X2 _26173_ (.A(_03087_),
    .B1(_03169_),
    .B2(_03171_),
    .C1(_03175_),
    .C2(_03075_),
    .ZN(_03176_));
 OR3_X2 _26174_ (.A1(_03165_),
    .A2(_03167_),
    .A3(_03176_),
    .ZN(_03177_));
 NAND4_X2 _26175_ (.A1(_03084_),
    .A2(_03125_),
    .A3(_03156_),
    .A4(_03177_),
    .ZN(_00120_));
 NAND2_X1 _26176_ (.A1(_03043_),
    .A2(_03029_),
    .ZN(_03178_));
 AOI21_X4 _26177_ (.A(net1037),
    .B1(_02981_),
    .B2(_02990_),
    .ZN(_03179_));
 NAND3_X1 _26178_ (.A1(_03072_),
    .A2(_03046_),
    .A3(_03047_),
    .ZN(_03180_));
 OAI21_X1 _26179_ (.A(_03180_),
    .B1(_02998_),
    .B2(_02972_),
    .ZN(_03181_));
 CLKBUF_X3 _26180_ (.A(_02974_),
    .Z(_03182_));
 AOI22_X1 _26181_ (.A1(_02976_),
    .A2(_03179_),
    .B1(_03181_),
    .B2(_03182_),
    .ZN(_03183_));
 OAI21_X4 _26182_ (.A(_03133_),
    .B1(_03049_),
    .B2(_03050_),
    .ZN(_03184_));
 INV_X2 _26183_ (.A(_15167_),
    .ZN(_03185_));
 OAI21_X1 _26184_ (.A(_03184_),
    .B1(_03070_),
    .B2(_03185_),
    .ZN(_03186_));
 AOI22_X2 _26185_ (.A1(_03072_),
    .A2(_03179_),
    .B1(_03186_),
    .B2(_03157_),
    .ZN(_03187_));
 NAND2_X2 _26186_ (.A1(_03015_),
    .A2(_03029_),
    .ZN(_03188_));
 AOI22_X1 _26187_ (.A1(net727),
    .A2(_03006_),
    .B1(_03111_),
    .B2(_03122_),
    .ZN(_03189_));
 NOR3_X4 _26188_ (.A1(_02968_),
    .A2(_02993_),
    .A3(_02996_),
    .ZN(_03190_));
 NOR2_X2 _26189_ (.A1(_03179_),
    .A2(_03190_),
    .ZN(_03191_));
 OAI21_X1 _26190_ (.A(_03189_),
    .B1(_03191_),
    .B2(_15169_),
    .ZN(_03192_));
 OAI222_X2 _26191_ (.A1(_03178_),
    .A2(_03183_),
    .B1(_03187_),
    .B2(_03188_),
    .C1(_03154_),
    .C2(_03192_),
    .ZN(_03193_));
 NAND2_X4 _26192_ (.A1(_03044_),
    .A2(_03032_),
    .ZN(_03194_));
 NAND2_X1 _26193_ (.A1(_03185_),
    .A2(_03117_),
    .ZN(_03195_));
 AOI21_X1 _26194_ (.A(_03182_),
    .B1(_03048_),
    .B2(_03195_),
    .ZN(_03196_));
 NAND3_X4 _26195_ (.A1(_03108_),
    .A2(_02982_),
    .A3(_02991_),
    .ZN(_03197_));
 AOI21_X4 _26196_ (.A(_02969_),
    .B1(_03197_),
    .B2(_03172_),
    .ZN(_03198_));
 NOR3_X1 _26197_ (.A1(_03194_),
    .A2(_03196_),
    .A3(_03198_),
    .ZN(_03199_));
 NOR3_X1 _26198_ (.A1(_03167_),
    .A2(_03193_),
    .A3(_03199_),
    .ZN(_03200_));
 AOI21_X1 _26199_ (.A(_03182_),
    .B1(_03048_),
    .B2(_03184_),
    .ZN(_03201_));
 AOI21_X1 _26200_ (.A(_03100_),
    .B1(_03117_),
    .B2(_03108_),
    .ZN(_03202_));
 OAI21_X1 _26201_ (.A(_03033_),
    .B1(_03202_),
    .B2(_03143_),
    .ZN(_03203_));
 AOI21_X4 _26202_ (.A(_03133_),
    .B1(_03046_),
    .B2(_03047_),
    .ZN(_03204_));
 NOR3_X4 _26203_ (.A1(_15176_),
    .A2(_02993_),
    .A3(_02996_),
    .ZN(_03205_));
 OAI21_X1 _26204_ (.A(_03157_),
    .B1(_03204_),
    .B2(_03205_),
    .ZN(_03206_));
 BUF_X8 _26205_ (.A(_03071_),
    .Z(_03207_));
 AOI21_X1 _26206_ (.A(_03100_),
    .B1(_03117_),
    .B2(_03207_),
    .ZN(_03208_));
 OAI21_X1 _26207_ (.A(_03206_),
    .B1(_03208_),
    .B2(_02975_),
    .ZN(_03209_));
 OAI22_X1 _26208_ (.A1(_03201_),
    .A2(_03203_),
    .B1(_03209_),
    .B2(_03194_),
    .ZN(_03210_));
 NOR2_X4 _26209_ (.A1(_03044_),
    .A2(_03086_),
    .ZN(_03211_));
 AOI21_X1 _26210_ (.A(_03037_),
    .B1(_03039_),
    .B2(_03207_),
    .ZN(_03212_));
 OAI221_X1 _26211_ (.A(_03211_),
    .B1(_03212_),
    .B2(_02970_),
    .C1(_03093_),
    .C2(_15169_),
    .ZN(_03213_));
 NOR3_X2 _26212_ (.A1(net1084),
    .A2(_03049_),
    .A3(_03050_),
    .ZN(_03214_));
 NOR3_X1 _26213_ (.A1(_03114_),
    .A2(_03214_),
    .A3(_03158_),
    .ZN(_03215_));
 INV_X1 _26214_ (.A(_03108_),
    .ZN(_03216_));
 NOR3_X1 _26215_ (.A1(_03216_),
    .A2(_03049_),
    .A3(_03050_),
    .ZN(_03217_));
 AOI21_X1 _26216_ (.A(_03217_),
    .B1(_03117_),
    .B2(_03000_),
    .ZN(_03218_));
 AOI21_X1 _26217_ (.A(_03215_),
    .B1(_03218_),
    .B2(_03143_),
    .ZN(_03219_));
 OAI21_X1 _26218_ (.A(_03213_),
    .B1(_03219_),
    .B2(_03188_),
    .ZN(_03220_));
 OAI21_X1 _26219_ (.A(_03060_),
    .B1(_03210_),
    .B2(_03220_),
    .ZN(_03221_));
 MUX2_X1 _26220_ (.A(_03094_),
    .B(_03207_),
    .S(_02973_),
    .Z(_03222_));
 NOR2_X2 _26221_ (.A1(_03222_),
    .A2(_03117_),
    .ZN(_03223_));
 NOR3_X1 _26222_ (.A1(_15186_),
    .A2(_02998_),
    .A3(_03086_),
    .ZN(_03224_));
 NOR3_X1 _26223_ (.A1(_03089_),
    .A2(_03223_),
    .A3(_03224_),
    .ZN(_03225_));
 OAI21_X1 _26224_ (.A(_02970_),
    .B1(_03099_),
    .B2(_03217_),
    .ZN(_03226_));
 MUX2_X1 _26225_ (.A(_03072_),
    .B(_02955_),
    .S(_02997_),
    .Z(_03227_));
 OAI21_X1 _26226_ (.A(_03226_),
    .B1(_03227_),
    .B2(_03143_),
    .ZN(_03228_));
 AOI21_X1 _26227_ (.A(_03225_),
    .B1(_03228_),
    .B2(_03033_),
    .ZN(_03229_));
 XNOR2_X1 _26228_ (.A(_02972_),
    .B(_02998_),
    .ZN(_03230_));
 AOI21_X1 _26229_ (.A(_03215_),
    .B1(_03230_),
    .B2(_03143_),
    .ZN(_03231_));
 AOI21_X1 _26230_ (.A(_03060_),
    .B1(_03231_),
    .B2(_03030_),
    .ZN(_03232_));
 AOI21_X2 _26231_ (.A(_03166_),
    .B1(_03232_),
    .B2(_03229_),
    .ZN(_03233_));
 CLKBUF_X3 _26232_ (.A(_03089_),
    .Z(_03234_));
 NOR3_X1 _26233_ (.A1(_03115_),
    .A2(_03037_),
    .A3(_03170_),
    .ZN(_03235_));
 AOI21_X1 _26234_ (.A(_03182_),
    .B1(_03116_),
    .B2(_03048_),
    .ZN(_03236_));
 NOR3_X1 _26235_ (.A1(_03076_),
    .A2(_03235_),
    .A3(_03236_),
    .ZN(_03237_));
 OAI21_X1 _26236_ (.A(_03032_),
    .B1(_02999_),
    .B2(_15190_),
    .ZN(_03238_));
 BUF_X4 _26237_ (.A(_03069_),
    .Z(_03239_));
 AOI21_X1 _26238_ (.A(_03239_),
    .B1(_03115_),
    .B2(_03185_),
    .ZN(_03240_));
 NAND2_X2 _26239_ (.A1(_02937_),
    .A2(_02973_),
    .ZN(_03241_));
 AOI21_X1 _26240_ (.A(_03238_),
    .B1(_03240_),
    .B2(_03241_),
    .ZN(_03242_));
 OAI21_X1 _26241_ (.A(_03234_),
    .B1(_03237_),
    .B2(_03242_),
    .ZN(_03243_));
 OAI21_X1 _26242_ (.A(_03115_),
    .B1(_03037_),
    .B2(_03170_),
    .ZN(_03244_));
 OAI21_X1 _26243_ (.A(_03244_),
    .B1(_03040_),
    .B2(_02971_),
    .ZN(_03245_));
 NOR2_X2 _26244_ (.A1(_03000_),
    .A2(_03117_),
    .ZN(_03246_));
 NOR2_X1 _26245_ (.A1(net515),
    .A2(_02998_),
    .ZN(_03247_));
 OAI21_X1 _26246_ (.A(_02971_),
    .B1(_03246_),
    .B2(_03247_),
    .ZN(_03248_));
 AOI21_X1 _26247_ (.A(_03076_),
    .B1(_03214_),
    .B2(_15159_),
    .ZN(_03249_));
 AOI22_X1 _26248_ (.A1(_03077_),
    .A2(_03245_),
    .B1(_03248_),
    .B2(_03249_),
    .ZN(_03250_));
 OAI21_X2 _26249_ (.A(_03243_),
    .B1(_03250_),
    .B2(_03234_),
    .ZN(_03251_));
 AOI221_X2 _26250_ (.A(_03200_),
    .B1(_03233_),
    .B2(_03221_),
    .C1(_03085_),
    .C2(_03251_),
    .ZN(_00121_));
 NOR3_X2 _26251_ (.A1(net563),
    .A2(_03049_),
    .A3(_03050_),
    .ZN(_03252_));
 NOR3_X1 _26252_ (.A1(_03092_),
    .A2(_03168_),
    .A3(_03252_),
    .ZN(_03253_));
 NOR3_X1 _26253_ (.A1(_03034_),
    .A2(_03158_),
    .A3(_03205_),
    .ZN(_03254_));
 OAI21_X1 _26254_ (.A(_03077_),
    .B1(_03253_),
    .B2(_03254_),
    .ZN(_03255_));
 AOI21_X1 _26255_ (.A(_15172_),
    .B1(_03046_),
    .B2(_03047_),
    .ZN(_03256_));
 NOR3_X1 _26256_ (.A1(_03092_),
    .A2(_03035_),
    .A3(_03256_),
    .ZN(_03257_));
 CLKBUF_X3 _26257_ (.A(_03239_),
    .Z(_03258_));
 AOI21_X1 _26258_ (.A(_03205_),
    .B1(_03258_),
    .B2(_15164_),
    .ZN(_03259_));
 AOI21_X1 _26259_ (.A(_03257_),
    .B1(_03259_),
    .B2(_15185_),
    .ZN(_03260_));
 OAI21_X1 _26260_ (.A(_03255_),
    .B1(_03260_),
    .B2(_03077_),
    .ZN(_03261_));
 NOR2_X1 _26261_ (.A1(_03097_),
    .A2(_03166_),
    .ZN(_03262_));
 NOR2_X1 _26262_ (.A1(_03097_),
    .A2(_03065_),
    .ZN(_03263_));
 NAND3_X1 _26263_ (.A1(_03143_),
    .A2(_03184_),
    .A3(_03197_),
    .ZN(_03264_));
 AOI21_X1 _26264_ (.A(_03144_),
    .B1(_02999_),
    .B2(_15164_),
    .ZN(_03265_));
 OAI21_X1 _26265_ (.A(_03264_),
    .B1(_03265_),
    .B2(_03092_),
    .ZN(_03266_));
 NOR2_X1 _26266_ (.A1(_02954_),
    .A2(_02968_),
    .ZN(_03267_));
 NOR3_X1 _26267_ (.A1(_02937_),
    .A2(_02997_),
    .A3(_03267_),
    .ZN(_03268_));
 NOR2_X1 _26268_ (.A1(net885),
    .A2(_02969_),
    .ZN(_03269_));
 MUX2_X1 _26269_ (.A(_02969_),
    .B(_02997_),
    .S(_02937_),
    .Z(_03270_));
 AOI221_X1 _26270_ (.A(_03268_),
    .B1(_03269_),
    .B2(_03116_),
    .C1(_03122_),
    .C2(_03270_),
    .ZN(_03271_));
 MUX2_X1 _26271_ (.A(_03266_),
    .B(_03271_),
    .S(_03088_),
    .Z(_03272_));
 AOI22_X1 _26272_ (.A1(_03261_),
    .A2(_03262_),
    .B1(_03263_),
    .B2(_03272_),
    .ZN(_03273_));
 AOI22_X1 _26273_ (.A1(_03046_),
    .A2(_03047_),
    .B1(_03029_),
    .B2(net725),
    .ZN(_03274_));
 OAI21_X1 _26274_ (.A(_03274_),
    .B1(_03086_),
    .B2(net727),
    .ZN(_03275_));
 OAI21_X1 _26275_ (.A(_03138_),
    .B1(_03086_),
    .B2(_03104_),
    .ZN(_03276_));
 OAI21_X1 _26276_ (.A(_03275_),
    .B1(_03276_),
    .B2(_03239_),
    .ZN(_03277_));
 AND3_X1 _26277_ (.A1(_03086_),
    .A2(_03184_),
    .A3(_03173_),
    .ZN(_03278_));
 OAI21_X1 _26278_ (.A(_02970_),
    .B1(_03087_),
    .B2(_03053_),
    .ZN(_03279_));
 OAI22_X2 _26279_ (.A1(_03092_),
    .A2(_03277_),
    .B1(_03278_),
    .B2(_03279_),
    .ZN(_03280_));
 NOR2_X1 _26280_ (.A1(_03089_),
    .A2(_03166_),
    .ZN(_03281_));
 NOR2_X1 _26281_ (.A1(_03090_),
    .A2(_03065_),
    .ZN(_03282_));
 AOI21_X1 _26282_ (.A(_03039_),
    .B1(_03087_),
    .B2(_03130_),
    .ZN(_03283_));
 MUX2_X1 _26283_ (.A(_03098_),
    .B(net727),
    .S(_03032_),
    .Z(_03284_));
 OAI221_X2 _26284_ (.A(_03283_),
    .B1(_03126_),
    .B2(_03087_),
    .C1(_03143_),
    .C2(_03284_),
    .ZN(_03285_));
 NAND2_X1 _26285_ (.A1(_15186_),
    .A2(_03032_),
    .ZN(_03286_));
 OAI21_X1 _26286_ (.A(_03286_),
    .B1(_03076_),
    .B2(_15183_),
    .ZN(_03287_));
 OAI21_X1 _26287_ (.A(_03285_),
    .B1(_03287_),
    .B2(_03258_),
    .ZN(_03288_));
 AOI221_X2 _26288_ (.A(_03141_),
    .B1(_03280_),
    .B2(_03281_),
    .C1(_03282_),
    .C2(_03288_),
    .ZN(_03289_));
 OAI21_X4 _26289_ (.A(_02975_),
    .B1(_03145_),
    .B2(_03006_),
    .ZN(_03290_));
 OAI21_X1 _26290_ (.A(_03143_),
    .B1(_02999_),
    .B2(_03080_),
    .ZN(_03291_));
 OAI211_X2 _26291_ (.A(_03090_),
    .B(_03290_),
    .C1(_03291_),
    .C2(_03246_),
    .ZN(_03292_));
 NOR2_X1 _26292_ (.A1(_02976_),
    .A2(_03054_),
    .ZN(_03293_));
 NAND3_X1 _26293_ (.A1(net516),
    .A2(_03046_),
    .A3(_03047_),
    .ZN(_03294_));
 OAI21_X1 _26294_ (.A(_03207_),
    .B1(_03049_),
    .B2(_03050_),
    .ZN(_03295_));
 AOI21_X1 _26295_ (.A(_03182_),
    .B1(_03294_),
    .B2(_03295_),
    .ZN(_03296_));
 OAI21_X1 _26296_ (.A(_03097_),
    .B1(_03293_),
    .B2(_03296_),
    .ZN(_03297_));
 AOI21_X1 _26297_ (.A(_03077_),
    .B1(_03292_),
    .B2(_03297_),
    .ZN(_03298_));
 MUX2_X1 _26298_ (.A(_03185_),
    .B(_15165_),
    .S(_02973_),
    .Z(_03299_));
 AOI21_X2 _26299_ (.A(_03044_),
    .B1(_03070_),
    .B2(_03299_),
    .ZN(_03300_));
 NAND2_X1 _26300_ (.A1(net725),
    .A2(_02969_),
    .ZN(_03301_));
 NAND3_X1 _26301_ (.A1(_02998_),
    .A2(_03301_),
    .A3(_03241_),
    .ZN(_03302_));
 NOR2_X1 _26302_ (.A1(_03099_),
    .A2(_03205_),
    .ZN(_03303_));
 AOI21_X1 _26303_ (.A(_03170_),
    .B1(_03069_),
    .B2(_02937_),
    .ZN(_03304_));
 MUX2_X1 _26304_ (.A(_03303_),
    .B(_03304_),
    .S(_02974_),
    .Z(_03305_));
 AOI221_X2 _26305_ (.A(_03087_),
    .B1(_03300_),
    .B2(_03302_),
    .C1(_03305_),
    .C2(_03089_),
    .ZN(_03306_));
 OR3_X2 _26306_ (.A1(_03166_),
    .A2(_03298_),
    .A3(_03306_),
    .ZN(_03307_));
 AOI22_X1 _26307_ (.A1(_15181_),
    .A2(_03121_),
    .B1(_03111_),
    .B2(net515),
    .ZN(_03308_));
 OAI21_X1 _26308_ (.A(_03166_),
    .B1(_03154_),
    .B2(_03308_),
    .ZN(_03309_));
 AOI21_X1 _26309_ (.A(_03188_),
    .B1(_03179_),
    .B2(_03053_),
    .ZN(_03310_));
 NAND3_X1 _26310_ (.A1(_15178_),
    .A2(_03184_),
    .A3(_03197_),
    .ZN(_03311_));
 AOI21_X1 _26311_ (.A(_03309_),
    .B1(_03310_),
    .B2(_03311_),
    .ZN(_03312_));
 NOR2_X1 _26312_ (.A1(_03098_),
    .A2(_02973_),
    .ZN(_03313_));
 NOR2_X1 _26313_ (.A1(_02998_),
    .A2(_03313_),
    .ZN(_03314_));
 AOI221_X1 _26314_ (.A(_03194_),
    .B1(_03241_),
    .B2(_03314_),
    .C1(_02999_),
    .C2(_15192_),
    .ZN(_03315_));
 CLKBUF_X3 _26315_ (.A(_03157_),
    .Z(_03316_));
 NOR2_X2 _26316_ (.A1(_03080_),
    .A2(_03053_),
    .ZN(_03317_));
 NAND3_X1 _26317_ (.A1(_03316_),
    .A2(_03258_),
    .A3(_03317_),
    .ZN(_03318_));
 INV_X1 _26318_ (.A(_03094_),
    .ZN(_03319_));
 OAI221_X1 _26319_ (.A(_03318_),
    .B1(_03191_),
    .B2(_03072_),
    .C1(_03319_),
    .C2(_03093_),
    .ZN(_03320_));
 AOI21_X1 _26320_ (.A(_03315_),
    .B1(_03320_),
    .B2(_03033_),
    .ZN(_03321_));
 AOI21_X1 _26321_ (.A(_03060_),
    .B1(_03312_),
    .B2(_03321_),
    .ZN(_03322_));
 AOI22_X2 _26322_ (.A1(_03273_),
    .A2(_03289_),
    .B1(_03307_),
    .B2(_03322_),
    .ZN(_00122_));
 NOR3_X4 _26323_ (.A1(_02974_),
    .A2(_02992_),
    .A3(_03035_),
    .ZN(_03323_));
 AOI21_X1 _26324_ (.A(_03162_),
    .B1(_03317_),
    .B2(_03117_),
    .ZN(_03324_));
 AOI21_X1 _26325_ (.A(_03323_),
    .B1(_03324_),
    .B2(_02975_),
    .ZN(_03325_));
 AOI22_X1 _26326_ (.A1(_15169_),
    .A2(_03190_),
    .B1(_03191_),
    .B2(net565),
    .ZN(_03326_));
 AOI221_X1 _26327_ (.A(_03142_),
    .B1(_03211_),
    .B2(_03325_),
    .C1(_03326_),
    .C2(_03045_),
    .ZN(_03327_));
 NAND3_X1 _26328_ (.A1(_15178_),
    .A2(_03079_),
    .A3(_03088_),
    .ZN(_03328_));
 NAND3_X1 _26329_ (.A1(_15185_),
    .A2(_03258_),
    .A3(_03077_),
    .ZN(_03329_));
 AOI21_X1 _26330_ (.A(_03122_),
    .B1(_03328_),
    .B2(_03329_),
    .ZN(_03330_));
 OR2_X1 _26331_ (.A1(_03094_),
    .A2(_03107_),
    .ZN(_03331_));
 NOR2_X2 _26332_ (.A1(_02937_),
    .A2(_03239_),
    .ZN(_03332_));
 AOI22_X1 _26333_ (.A1(net1045),
    .A2(_03258_),
    .B1(_03332_),
    .B2(_03076_),
    .ZN(_03333_));
 OAI221_X1 _26334_ (.A(_03234_),
    .B1(_03093_),
    .B2(_03331_),
    .C1(_03333_),
    .C2(_15185_),
    .ZN(_03334_));
 OAI21_X1 _26335_ (.A(_03327_),
    .B1(_03330_),
    .B2(_03334_),
    .ZN(_03335_));
 NOR2_X2 _26336_ (.A1(_03141_),
    .A2(_03065_),
    .ZN(_03336_));
 AOI221_X1 _26337_ (.A(_03032_),
    .B1(_03111_),
    .B2(_03094_),
    .C1(_15159_),
    .C2(_03168_),
    .ZN(_03337_));
 NAND3_X1 _26338_ (.A1(_03234_),
    .A2(_03290_),
    .A3(_03337_),
    .ZN(_03338_));
 NOR3_X1 _26339_ (.A1(_03034_),
    .A2(_02992_),
    .A3(_03252_),
    .ZN(_03339_));
 AOI21_X2 _26340_ (.A(_03145_),
    .B1(_03239_),
    .B2(_03000_),
    .ZN(_03340_));
 AOI21_X2 _26341_ (.A(_03339_),
    .B1(_03340_),
    .B2(_15178_),
    .ZN(_03341_));
 OAI21_X1 _26342_ (.A(_03338_),
    .B1(_03341_),
    .B2(_03194_),
    .ZN(_03342_));
 OAI21_X1 _26343_ (.A(_15185_),
    .B1(_03099_),
    .B2(_03162_),
    .ZN(_03343_));
 OR3_X1 _26344_ (.A1(_02971_),
    .A2(_03144_),
    .A3(_03147_),
    .ZN(_03344_));
 NAND3_X1 _26345_ (.A1(_03045_),
    .A2(_03343_),
    .A3(_03344_),
    .ZN(_03345_));
 AOI21_X1 _26346_ (.A(_03267_),
    .B1(_15158_),
    .B2(_15164_),
    .ZN(_03346_));
 OAI221_X1 _26347_ (.A(_03211_),
    .B1(_03346_),
    .B2(_03258_),
    .C1(_03102_),
    .C2(_03098_),
    .ZN(_03347_));
 NAND2_X1 _26348_ (.A1(_03345_),
    .A2(_03347_),
    .ZN(_03348_));
 OAI21_X2 _26349_ (.A(_03336_),
    .B1(_03348_),
    .B2(_03342_),
    .ZN(_03349_));
 NOR2_X1 _26350_ (.A1(_03079_),
    .A2(_03138_),
    .ZN(_03350_));
 INV_X1 _26351_ (.A(_02976_),
    .ZN(_03351_));
 NAND3_X2 _26352_ (.A1(_03351_),
    .A2(_03046_),
    .A3(_03047_),
    .ZN(_03352_));
 NAND2_X1 _26353_ (.A1(_15185_),
    .A2(_03352_),
    .ZN(_03353_));
 NAND3_X4 _26354_ (.A1(_03036_),
    .A2(_02982_),
    .A3(_02991_),
    .ZN(_03354_));
 OAI21_X4 _26355_ (.A(_15172_),
    .B1(_03003_),
    .B2(_03004_),
    .ZN(_03355_));
 AND2_X2 _26356_ (.A1(_03354_),
    .A2(_03355_),
    .ZN(_03356_));
 MUX2_X1 _26357_ (.A(_03035_),
    .B(_03356_),
    .S(_03107_),
    .Z(_03357_));
 OAI221_X2 _26358_ (.A(_03234_),
    .B1(_03350_),
    .B2(_03353_),
    .C1(_03357_),
    .C2(_15185_),
    .ZN(_03358_));
 AND2_X1 _26359_ (.A1(_02974_),
    .A2(_03317_),
    .ZN(_03359_));
 OAI21_X1 _26360_ (.A(_03258_),
    .B1(_03034_),
    .B2(net565),
    .ZN(_03360_));
 OAI221_X1 _26361_ (.A(_03211_),
    .B1(_03359_),
    .B2(_03360_),
    .C1(_03222_),
    .C2(_03258_),
    .ZN(_03361_));
 AOI21_X1 _26362_ (.A(_03188_),
    .B1(_03111_),
    .B2(_15164_),
    .ZN(_03362_));
 NOR2_X1 _26363_ (.A1(_03092_),
    .A2(_03332_),
    .ZN(_03363_));
 OAI221_X1 _26364_ (.A(_03362_),
    .B1(_03363_),
    .B2(_15158_),
    .C1(_03108_),
    .C2(_03054_),
    .ZN(_03364_));
 NAND4_X2 _26365_ (.A1(_03067_),
    .A2(_03358_),
    .A3(_03361_),
    .A4(_03364_),
    .ZN(_03365_));
 AOI21_X1 _26366_ (.A(_03037_),
    .B1(_03079_),
    .B2(_15159_),
    .ZN(_03366_));
 OAI221_X1 _26367_ (.A(_03030_),
    .B1(_03151_),
    .B2(_15169_),
    .C1(_03366_),
    .C2(_15178_),
    .ZN(_03367_));
 AOI21_X2 _26368_ (.A(_03134_),
    .B1(_03046_),
    .B2(_03047_),
    .ZN(_03368_));
 AOI222_X2 _26369_ (.A1(_03122_),
    .A2(_03368_),
    .B1(_03078_),
    .B2(_03048_),
    .C1(_03127_),
    .C2(_03332_),
    .ZN(_03369_));
 OAI21_X1 _26370_ (.A(_03367_),
    .B1(_03369_),
    .B2(_03154_),
    .ZN(_03370_));
 NOR3_X1 _26371_ (.A1(_03094_),
    .A2(_03049_),
    .A3(_03050_),
    .ZN(_03371_));
 OAI21_X1 _26372_ (.A(_02975_),
    .B1(_03109_),
    .B2(_03371_),
    .ZN(_03372_));
 NAND3_X1 _26373_ (.A1(_02971_),
    .A2(_03048_),
    .A3(_03172_),
    .ZN(_03373_));
 AND3_X1 _26374_ (.A1(_03090_),
    .A2(_03372_),
    .A3(_03373_),
    .ZN(_03374_));
 NOR3_X1 _26375_ (.A1(_02971_),
    .A2(_02992_),
    .A3(_03145_),
    .ZN(_03375_));
 AOI211_X2 _26376_ (.A(_02974_),
    .B(_03158_),
    .C1(_03039_),
    .C2(_03000_),
    .ZN(_03376_));
 NOR3_X1 _26377_ (.A1(_03375_),
    .A2(_03234_),
    .A3(_03376_),
    .ZN(_03377_));
 NOR3_X1 _26378_ (.A1(_03077_),
    .A2(_03374_),
    .A3(_03377_),
    .ZN(_03378_));
 OAI21_X1 _26379_ (.A(_03085_),
    .B1(_03370_),
    .B2(_03378_),
    .ZN(_03379_));
 NAND4_X2 _26380_ (.A1(_03379_),
    .A2(_03349_),
    .A3(_03365_),
    .A4(_03335_),
    .ZN(_00123_));
 AOI21_X1 _26381_ (.A(_03076_),
    .B1(_03034_),
    .B2(_03104_),
    .ZN(_03380_));
 AOI21_X1 _26382_ (.A(_03097_),
    .B1(_03244_),
    .B2(_03380_),
    .ZN(_03381_));
 OAI21_X1 _26383_ (.A(_15178_),
    .B1(_03099_),
    .B2(_03170_),
    .ZN(_03382_));
 AOI21_X1 _26384_ (.A(_03205_),
    .B1(_03239_),
    .B2(_03000_),
    .ZN(_03383_));
 OAI21_X1 _26385_ (.A(_03382_),
    .B1(_03383_),
    .B2(_15178_),
    .ZN(_03384_));
 OAI21_X1 _26386_ (.A(_03381_),
    .B1(_03384_),
    .B2(_03088_),
    .ZN(_03385_));
 AOI21_X1 _26387_ (.A(_03143_),
    .B1(_03051_),
    .B2(_03352_),
    .ZN(_03386_));
 AOI21_X1 _26388_ (.A(_03386_),
    .B1(_03356_),
    .B2(_03092_),
    .ZN(_03387_));
 OR2_X1 _26389_ (.A1(_03188_),
    .A2(_03387_),
    .ZN(_03388_));
 AOI21_X1 _26390_ (.A(_03088_),
    .B1(_03078_),
    .B2(_03258_),
    .ZN(_03389_));
 NAND2_X1 _26391_ (.A1(_03113_),
    .A2(_03389_),
    .ZN(_03390_));
 NAND4_X1 _26392_ (.A1(_03085_),
    .A2(_03385_),
    .A3(_03388_),
    .A4(_03390_),
    .ZN(_03391_));
 AOI21_X1 _26393_ (.A(_03005_),
    .B1(_03239_),
    .B2(_15164_),
    .ZN(_03392_));
 OAI221_X1 _26394_ (.A(_03089_),
    .B1(_03102_),
    .B2(_03104_),
    .C1(_03392_),
    .C2(_02971_),
    .ZN(_03393_));
 MUX2_X1 _26395_ (.A(_03072_),
    .B(_03301_),
    .S(_03239_),
    .Z(_03394_));
 OAI21_X1 _26396_ (.A(_03393_),
    .B1(_03394_),
    .B2(_03090_),
    .ZN(_03395_));
 NAND2_X1 _26397_ (.A1(_03116_),
    .A2(_03197_),
    .ZN(_03396_));
 AOI221_X1 _26398_ (.A(_03044_),
    .B1(_03190_),
    .B2(_03118_),
    .C1(_03396_),
    .C2(_03134_),
    .ZN(_03397_));
 OAI22_X2 _26399_ (.A1(net1084),
    .A2(_03054_),
    .B1(_03093_),
    .B2(_02937_),
    .ZN(_03398_));
 OAI21_X1 _26400_ (.A(_03116_),
    .B1(_02974_),
    .B2(_02937_),
    .ZN(_03399_));
 AOI211_X2 _26401_ (.A(_03015_),
    .B(_03398_),
    .C1(_03399_),
    .C2(_03104_),
    .ZN(_03400_));
 NAND2_X1 _26402_ (.A1(_03043_),
    .A2(_03069_),
    .ZN(_03401_));
 NAND3_X1 _26403_ (.A1(_03080_),
    .A2(_03096_),
    .A3(_03039_),
    .ZN(_03402_));
 AOI21_X1 _26404_ (.A(_02971_),
    .B1(_03401_),
    .B2(_03402_),
    .ZN(_03403_));
 NAND4_X1 _26405_ (.A1(_03216_),
    .A2(_02970_),
    .A3(_03096_),
    .A4(_03039_),
    .ZN(_03404_));
 OR2_X1 _26406_ (.A1(_03096_),
    .A2(_03355_),
    .ZN(_03405_));
 OAI21_X1 _26407_ (.A(_03000_),
    .B1(_03157_),
    .B2(_03096_),
    .ZN(_03406_));
 NAND4_X1 _26408_ (.A1(_15158_),
    .A2(_03404_),
    .A3(_03405_),
    .A4(_03406_),
    .ZN(_03407_));
 OAI22_X1 _26409_ (.A1(_03397_),
    .A2(_03400_),
    .B1(_03403_),
    .B2(_03407_),
    .ZN(_03408_));
 MUX2_X1 _26410_ (.A(_03395_),
    .B(_03408_),
    .S(_03077_),
    .Z(_03409_));
 NAND2_X1 _26411_ (.A1(_03134_),
    .A2(_03044_),
    .ZN(_03410_));
 OAI221_X1 _26412_ (.A(_03239_),
    .B1(_03241_),
    .B2(_03044_),
    .C1(_03410_),
    .C2(_03216_),
    .ZN(_03411_));
 AOI21_X1 _26413_ (.A(_15169_),
    .B1(_03134_),
    .B2(_03096_),
    .ZN(_03412_));
 OAI21_X1 _26414_ (.A(_03127_),
    .B1(_03412_),
    .B2(_03000_),
    .ZN(_03413_));
 OAI21_X1 _26415_ (.A(_03411_),
    .B1(_03413_),
    .B2(_03121_),
    .ZN(_03414_));
 OAI21_X1 _26416_ (.A(_03169_),
    .B1(_03096_),
    .B2(_02970_),
    .ZN(_03415_));
 AOI21_X1 _26417_ (.A(_03087_),
    .B1(_03415_),
    .B2(_15159_),
    .ZN(_03416_));
 OAI21_X1 _26418_ (.A(_03197_),
    .B1(_02998_),
    .B2(net727),
    .ZN(_03417_));
 OAI21_X1 _26419_ (.A(_03127_),
    .B1(_03417_),
    .B2(_03182_),
    .ZN(_03418_));
 OAI21_X1 _26420_ (.A(_03355_),
    .B1(_03100_),
    .B2(_02970_),
    .ZN(_03419_));
 MUX2_X1 _26421_ (.A(_03418_),
    .B(_03419_),
    .S(_03089_),
    .Z(_03420_));
 AOI221_X1 _26422_ (.A(_03065_),
    .B1(_03414_),
    .B2(_03416_),
    .C1(_03420_),
    .C2(_03088_),
    .ZN(_03421_));
 AOI22_X1 _26423_ (.A1(_15158_),
    .A2(_03190_),
    .B1(_03352_),
    .B2(_03092_),
    .ZN(_03422_));
 OAI21_X1 _26424_ (.A(_03065_),
    .B1(_03154_),
    .B2(_03422_),
    .ZN(_03423_));
 NOR2_X1 _26425_ (.A1(_03185_),
    .A2(_02970_),
    .ZN(_03424_));
 OAI21_X1 _26426_ (.A(_02999_),
    .B1(_03130_),
    .B2(_03424_),
    .ZN(_03425_));
 AND2_X1 _26427_ (.A1(_03074_),
    .A2(_03425_),
    .ZN(_03426_));
 NOR2_X1 _26428_ (.A1(_03208_),
    .A2(_03410_),
    .ZN(_03427_));
 MUX2_X1 _26429_ (.A(_03053_),
    .B(_03216_),
    .S(_03039_),
    .Z(_03428_));
 NOR2_X1 _26430_ (.A1(_03092_),
    .A2(_03428_),
    .ZN(_03429_));
 NOR2_X1 _26431_ (.A1(_02975_),
    .A2(_03230_),
    .ZN(_03430_));
 OAI33_X1 _26432_ (.A1(_03077_),
    .A2(_03426_),
    .A3(_03427_),
    .B1(_03429_),
    .B2(_03430_),
    .B3(_03194_),
    .ZN(_03431_));
 OAI21_X1 _26433_ (.A(_03060_),
    .B1(_03423_),
    .B2(_03431_),
    .ZN(_03432_));
 OAI221_X1 _26434_ (.A(_03391_),
    .B1(_03409_),
    .B2(_03142_),
    .C1(_03421_),
    .C2(_03432_),
    .ZN(_00124_));
 AOI21_X2 _26435_ (.A(_03144_),
    .B1(_02997_),
    .B2(_02976_),
    .ZN(_03433_));
 OAI221_X2 _26436_ (.A(_03089_),
    .B1(_03151_),
    .B2(_03207_),
    .C1(_03433_),
    .C2(_03157_),
    .ZN(_03434_));
 MUX2_X1 _26437_ (.A(_03071_),
    .B(_02954_),
    .S(_02968_),
    .Z(_03435_));
 NOR2_X1 _26438_ (.A1(_03043_),
    .A2(_02997_),
    .ZN(_03436_));
 NOR2_X1 _26439_ (.A1(_03185_),
    .A2(net1037),
    .ZN(_03437_));
 NOR3_X2 _26440_ (.A1(_03043_),
    .A2(_03068_),
    .A3(_03437_),
    .ZN(_03438_));
 AOI221_X2 _26441_ (.A(_03029_),
    .B1(_03435_),
    .B2(_03436_),
    .C1(_03438_),
    .C2(_03127_),
    .ZN(_03439_));
 OAI22_X1 _26442_ (.A1(_15159_),
    .A2(_03048_),
    .B1(_03190_),
    .B2(_15158_),
    .ZN(_03440_));
 AOI221_X2 _26443_ (.A(_03066_),
    .B1(_03434_),
    .B2(_03439_),
    .C1(_03440_),
    .C2(_03045_),
    .ZN(_03441_));
 AOI22_X1 _26444_ (.A1(_03053_),
    .A2(_02998_),
    .B1(_03051_),
    .B2(_03114_),
    .ZN(_03442_));
 OAI21_X1 _26445_ (.A(_03336_),
    .B1(_03442_),
    .B2(_03194_),
    .ZN(_03443_));
 NAND2_X1 _26446_ (.A1(_03182_),
    .A2(_03356_),
    .ZN(_03444_));
 AOI21_X1 _26447_ (.A(_03154_),
    .B1(_03006_),
    .B2(_03134_),
    .ZN(_03445_));
 MUX2_X1 _26448_ (.A(_03351_),
    .B(_02937_),
    .S(_02997_),
    .Z(_03446_));
 AOI21_X1 _26449_ (.A(_03188_),
    .B1(_03446_),
    .B2(_03115_),
    .ZN(_03447_));
 AOI221_X2 _26450_ (.A(_03443_),
    .B1(_03444_),
    .B2(_03445_),
    .C1(_03447_),
    .C2(_03159_),
    .ZN(_03448_));
 OAI21_X1 _26451_ (.A(_03178_),
    .B1(_03441_),
    .B2(_03448_),
    .ZN(_03449_));
 MUX2_X1 _26452_ (.A(_03094_),
    .B(_03359_),
    .S(_03086_),
    .Z(_03450_));
 NOR2_X1 _26453_ (.A1(_03079_),
    .A2(_03450_),
    .ZN(_03451_));
 AOI221_X1 _26454_ (.A(_03117_),
    .B1(_03086_),
    .B2(_03313_),
    .C1(_03157_),
    .C2(_03207_),
    .ZN(_03452_));
 NOR3_X1 _26455_ (.A1(_03234_),
    .A2(_03451_),
    .A3(_03452_),
    .ZN(_03453_));
 OAI22_X2 _26456_ (.A1(_02976_),
    .A2(_03102_),
    .B1(_03437_),
    .B2(_03121_),
    .ZN(_03454_));
 AOI21_X1 _26457_ (.A(_03166_),
    .B1(_03454_),
    .B2(_03033_),
    .ZN(_03455_));
 NAND3_X1 _26458_ (.A1(_03316_),
    .A2(_03184_),
    .A3(_03354_),
    .ZN(_03456_));
 OAI21_X1 _26459_ (.A(_03456_),
    .B1(_03433_),
    .B2(_03034_),
    .ZN(_03457_));
 OAI21_X1 _26460_ (.A(_03455_),
    .B1(_03457_),
    .B2(_03194_),
    .ZN(_03458_));
 AOI21_X1 _26461_ (.A(_15158_),
    .B1(_03096_),
    .B2(_15159_),
    .ZN(_03459_));
 OAI221_X2 _26462_ (.A(_03107_),
    .B1(_03401_),
    .B2(_03222_),
    .C1(_03459_),
    .C2(_03093_),
    .ZN(_03460_));
 XNOR2_X1 _26463_ (.A(_03090_),
    .B(_03214_),
    .ZN(_03461_));
 AOI21_X1 _26464_ (.A(_03460_),
    .B1(_03461_),
    .B2(_15164_),
    .ZN(_03462_));
 AOI21_X1 _26465_ (.A(_03204_),
    .B1(_02999_),
    .B2(net1045),
    .ZN(_03463_));
 OAI221_X1 _26466_ (.A(_03030_),
    .B1(_03151_),
    .B2(_15164_),
    .C1(_03463_),
    .C2(_03034_),
    .ZN(_03464_));
 AOI21_X1 _26467_ (.A(_03109_),
    .B1(_02999_),
    .B2(_02976_),
    .ZN(_03465_));
 OAI221_X1 _26468_ (.A(_03211_),
    .B1(_03465_),
    .B2(_03316_),
    .C1(_03054_),
    .C2(_03122_),
    .ZN(_03466_));
 NAND3_X1 _26469_ (.A1(_03166_),
    .A2(_03464_),
    .A3(_03466_),
    .ZN(_03467_));
 OAI221_X1 _26470_ (.A(_03141_),
    .B1(_03453_),
    .B2(_03458_),
    .C1(_03467_),
    .C2(_03462_),
    .ZN(_03468_));
 OAI21_X1 _26471_ (.A(_15185_),
    .B1(_03099_),
    .B2(_03252_),
    .ZN(_03469_));
 OAI21_X1 _26472_ (.A(_03469_),
    .B1(_03366_),
    .B2(_15185_),
    .ZN(_03470_));
 NOR2_X1 _26473_ (.A1(_03115_),
    .A2(_03091_),
    .ZN(_03471_));
 AOI221_X1 _26474_ (.A(_03471_),
    .B1(_03111_),
    .B2(net565),
    .C1(_03258_),
    .C2(_03053_),
    .ZN(_03472_));
 AOI22_X1 _26475_ (.A1(_03441_),
    .A2(_03470_),
    .B1(_03472_),
    .B2(_03448_),
    .ZN(_03473_));
 AND3_X2 _26476_ (.A1(_03449_),
    .A2(_03468_),
    .A3(_03473_),
    .ZN(_00125_));
 NOR2_X1 _26477_ (.A1(_03122_),
    .A2(_03115_),
    .ZN(_03474_));
 OR2_X1 _26478_ (.A1(_03117_),
    .A2(_03313_),
    .ZN(_03475_));
 OAI221_X1 _26479_ (.A(_03107_),
    .B1(_03474_),
    .B2(_03475_),
    .C1(_03079_),
    .C2(_15181_),
    .ZN(_03476_));
 AOI21_X1 _26480_ (.A(_03371_),
    .B1(_03121_),
    .B2(_15159_),
    .ZN(_03477_));
 OAI221_X1 _26481_ (.A(_03076_),
    .B1(_03054_),
    .B2(net515),
    .C1(_03477_),
    .C2(_03316_),
    .ZN(_03478_));
 NAND3_X1 _26482_ (.A1(_03476_),
    .A2(_03234_),
    .A3(_03478_),
    .ZN(_03479_));
 AOI21_X1 _26483_ (.A(_03182_),
    .B1(_03116_),
    .B2(_03354_),
    .ZN(_03480_));
 NOR2_X1 _26484_ (.A1(_03070_),
    .A2(_03317_),
    .ZN(_03481_));
 NOR3_X1 _26485_ (.A1(_03115_),
    .A2(_03247_),
    .A3(_03481_),
    .ZN(_03482_));
 OR3_X1 _26486_ (.A1(_03154_),
    .A2(_03480_),
    .A3(_03482_),
    .ZN(_03483_));
 AND2_X1 _26487_ (.A1(_03316_),
    .A2(_03340_),
    .ZN(_03484_));
 NOR2_X1 _26488_ (.A1(_03316_),
    .A2(_03101_),
    .ZN(_03485_));
 OAI21_X1 _26489_ (.A(_03045_),
    .B1(_03484_),
    .B2(_03485_),
    .ZN(_03486_));
 AND4_X2 _26490_ (.A1(_03085_),
    .A2(_03479_),
    .A3(_03483_),
    .A4(_03486_),
    .ZN(_03487_));
 AOI21_X1 _26491_ (.A(_03256_),
    .B1(_03079_),
    .B2(_03094_),
    .ZN(_03488_));
 OAI221_X1 _26492_ (.A(_03090_),
    .B1(_03054_),
    .B2(_15164_),
    .C1(_03488_),
    .C2(_15178_),
    .ZN(_03489_));
 NOR2_X1 _26493_ (.A1(_03088_),
    .A2(_03300_),
    .ZN(_03490_));
 NAND2_X1 _26494_ (.A1(_03489_),
    .A2(_03490_),
    .ZN(_03491_));
 OAI21_X1 _26495_ (.A(_03090_),
    .B1(_03150_),
    .B2(_03323_),
    .ZN(_03492_));
 AOI21_X1 _26496_ (.A(_03089_),
    .B1(_03121_),
    .B2(_15180_),
    .ZN(_03493_));
 OAI21_X1 _26497_ (.A(_03079_),
    .B1(_03316_),
    .B2(_03104_),
    .ZN(_03494_));
 OAI21_X1 _26498_ (.A(_03493_),
    .B1(_03494_),
    .B2(_03269_),
    .ZN(_03495_));
 NAND3_X1 _26499_ (.A1(_03088_),
    .A2(_03492_),
    .A3(_03495_),
    .ZN(_03496_));
 AOI21_X1 _26500_ (.A(_03142_),
    .B1(_03491_),
    .B2(_03496_),
    .ZN(_03497_));
 OAI21_X1 _26501_ (.A(_03355_),
    .B1(_03070_),
    .B2(_03108_),
    .ZN(_03498_));
 AOI221_X2 _26502_ (.A(_03032_),
    .B1(_03179_),
    .B2(net1045),
    .C1(_03498_),
    .C2(_03157_),
    .ZN(_03499_));
 NAND3_X1 _26503_ (.A1(_03316_),
    .A2(_03048_),
    .A3(_03355_),
    .ZN(_03500_));
 OAI22_X2 _26504_ (.A1(_03080_),
    .A2(_03053_),
    .B1(_03049_),
    .B2(_03050_),
    .ZN(_03501_));
 OAI21_X1 _26505_ (.A(_03501_),
    .B1(_03121_),
    .B2(_03122_),
    .ZN(_03502_));
 OAI21_X1 _26506_ (.A(_03500_),
    .B1(_03502_),
    .B2(_03034_),
    .ZN(_03503_));
 AOI21_X1 _26507_ (.A(_03499_),
    .B1(_03503_),
    .B2(_03077_),
    .ZN(_03504_));
 NAND2_X1 _26508_ (.A1(_03234_),
    .A2(_03336_),
    .ZN(_03505_));
 NAND2_X1 _26509_ (.A1(_03097_),
    .A2(_03336_),
    .ZN(_03506_));
 AOI21_X1 _26510_ (.A(_03205_),
    .B1(_03070_),
    .B2(_03118_),
    .ZN(_03507_));
 OAI21_X1 _26511_ (.A(_03173_),
    .B1(_02998_),
    .B2(_03207_),
    .ZN(_03508_));
 MUX2_X1 _26512_ (.A(_03507_),
    .B(_03508_),
    .S(_03134_),
    .Z(_03509_));
 NOR3_X1 _26513_ (.A1(_15179_),
    .A2(_15188_),
    .A3(_03070_),
    .ZN(_03510_));
 MUX2_X1 _26514_ (.A(net1084),
    .B(_03114_),
    .S(_02972_),
    .Z(_03511_));
 AOI21_X1 _26515_ (.A(_03510_),
    .B1(_03511_),
    .B2(_03239_),
    .ZN(_03512_));
 MUX2_X1 _26516_ (.A(_03509_),
    .B(_03512_),
    .S(_03107_),
    .Z(_03513_));
 OAI22_X2 _26517_ (.A1(_03504_),
    .A2(_03505_),
    .B1(_03506_),
    .B2(_03513_),
    .ZN(_03514_));
 OAI21_X1 _26518_ (.A(_15164_),
    .B1(_03316_),
    .B2(_03168_),
    .ZN(_03515_));
 AOI22_X1 _26519_ (.A1(_15169_),
    .A2(_03368_),
    .B1(_03111_),
    .B2(net516),
    .ZN(_03516_));
 NAND3_X1 _26520_ (.A1(_03107_),
    .A2(_03515_),
    .A3(_03516_),
    .ZN(_03517_));
 AND3_X1 _26521_ (.A1(_03157_),
    .A2(_03354_),
    .A3(_03355_),
    .ZN(_03518_));
 NOR2_X1 _26522_ (.A1(_03182_),
    .A2(_03168_),
    .ZN(_03519_));
 OR3_X1 _26523_ (.A1(_03087_),
    .A2(_03518_),
    .A3(_03519_),
    .ZN(_03520_));
 NAND3_X1 _26524_ (.A1(_03097_),
    .A2(_03517_),
    .A3(_03520_),
    .ZN(_03521_));
 AOI21_X1 _26525_ (.A(_03267_),
    .B1(_03114_),
    .B2(_03098_),
    .ZN(_03522_));
 MUX2_X1 _26526_ (.A(_15190_),
    .B(_03522_),
    .S(_03039_),
    .Z(_03523_));
 OAI21_X1 _26527_ (.A(_03107_),
    .B1(_03126_),
    .B2(_03079_),
    .ZN(_03524_));
 OAI22_X1 _26528_ (.A1(_15158_),
    .A2(_03316_),
    .B1(_03151_),
    .B2(_02976_),
    .ZN(_03525_));
 OAI221_X1 _26529_ (.A(_03234_),
    .B1(_03088_),
    .B2(_03523_),
    .C1(_03524_),
    .C2(_03525_),
    .ZN(_03526_));
 AOI21_X1 _26530_ (.A(_03066_),
    .B1(_03521_),
    .B2(_03526_),
    .ZN(_03527_));
 NOR4_X4 _26531_ (.A1(_03527_),
    .A2(_03497_),
    .A3(_03514_),
    .A4(_03487_),
    .ZN(_00126_));
 OAI21_X1 _26532_ (.A(_03354_),
    .B1(_03401_),
    .B2(_03098_),
    .ZN(_03528_));
 NAND2_X1 _26533_ (.A1(_03182_),
    .A2(_03528_),
    .ZN(_03529_));
 OAI21_X1 _26534_ (.A(_03093_),
    .B1(_02997_),
    .B2(_03043_),
    .ZN(_03530_));
 AOI221_X2 _26535_ (.A(_03029_),
    .B1(_03530_),
    .B2(_03207_),
    .C1(_02969_),
    .C2(_03014_),
    .ZN(_03531_));
 NOR4_X1 _26536_ (.A1(_03207_),
    .A2(_02973_),
    .A3(_03043_),
    .A4(_03069_),
    .ZN(_03532_));
 NOR2_X1 _26537_ (.A1(_15169_),
    .A2(_03114_),
    .ZN(_03533_));
 AOI21_X1 _26538_ (.A(_03532_),
    .B1(_03533_),
    .B2(_03129_),
    .ZN(_03534_));
 NOR2_X1 _26539_ (.A1(_03015_),
    .A2(_03069_),
    .ZN(_03535_));
 AOI21_X1 _26540_ (.A(_03535_),
    .B1(_03436_),
    .B2(net727),
    .ZN(_03536_));
 NOR3_X1 _26541_ (.A1(_03114_),
    .A2(_03043_),
    .A3(_03069_),
    .ZN(_03537_));
 NOR2_X1 _26542_ (.A1(_03179_),
    .A2(_03537_),
    .ZN(_03538_));
 OAI221_X2 _26543_ (.A(_03534_),
    .B1(_03536_),
    .B2(_15158_),
    .C1(_03538_),
    .C2(_03000_),
    .ZN(_03539_));
 AOI221_X2 _26544_ (.A(_03142_),
    .B1(_03529_),
    .B2(_03531_),
    .C1(_03539_),
    .C2(_03087_),
    .ZN(_03540_));
 AOI21_X1 _26545_ (.A(_03143_),
    .B1(_03294_),
    .B2(_03195_),
    .ZN(_03541_));
 OAI21_X1 _26546_ (.A(_03090_),
    .B1(_03430_),
    .B2(_03541_),
    .ZN(_03542_));
 OAI221_X1 _26547_ (.A(_03097_),
    .B1(_03079_),
    .B2(_03207_),
    .C1(_03093_),
    .C2(_03118_),
    .ZN(_03543_));
 NAND3_X1 _26548_ (.A1(_03088_),
    .A2(_03542_),
    .A3(_03543_),
    .ZN(_03544_));
 NOR2_X1 _26549_ (.A1(_03104_),
    .A2(_03134_),
    .ZN(_03545_));
 NOR3_X1 _26550_ (.A1(_03121_),
    .A2(_03130_),
    .A3(_03545_),
    .ZN(_03546_));
 OAI21_X1 _26551_ (.A(_03211_),
    .B1(_02999_),
    .B2(_15188_),
    .ZN(_03547_));
 OAI21_X1 _26552_ (.A(_03085_),
    .B1(_03546_),
    .B2(_03547_),
    .ZN(_03548_));
 NOR2_X1 _26553_ (.A1(_03246_),
    .A2(_03037_),
    .ZN(_03549_));
 AOI21_X1 _26554_ (.A(_03201_),
    .B1(_03549_),
    .B2(_03034_),
    .ZN(_03550_));
 AOI21_X1 _26555_ (.A(_03548_),
    .B1(_03550_),
    .B2(_03030_),
    .ZN(_03551_));
 NOR2_X1 _26556_ (.A1(_03108_),
    .A2(_02969_),
    .ZN(_03552_));
 AOI21_X1 _26557_ (.A(_03100_),
    .B1(_03069_),
    .B2(_02937_),
    .ZN(_03553_));
 AOI21_X1 _26558_ (.A(_03552_),
    .B1(_03553_),
    .B2(_03114_),
    .ZN(_03554_));
 NOR3_X1 _26559_ (.A1(_02974_),
    .A2(_03144_),
    .A3(_03147_),
    .ZN(_03555_));
 OR2_X2 _26560_ (.A1(_03198_),
    .A2(_03555_),
    .ZN(_03556_));
 AOI221_X2 _26561_ (.A(_03065_),
    .B1(_03211_),
    .B2(_03554_),
    .C1(_03045_),
    .C2(_03556_),
    .ZN(_03557_));
 OAI21_X1 _26562_ (.A(_03501_),
    .B1(_03070_),
    .B2(_02937_),
    .ZN(_03558_));
 NAND2_X1 _26563_ (.A1(_03180_),
    .A2(_03355_),
    .ZN(_03559_));
 MUX2_X1 _26564_ (.A(_03558_),
    .B(_03559_),
    .S(_03134_),
    .Z(_03560_));
 AOI21_X1 _26565_ (.A(_03170_),
    .B1(_03511_),
    .B2(_03121_),
    .ZN(_03561_));
 MUX2_X1 _26566_ (.A(_03560_),
    .B(_03561_),
    .S(_03076_),
    .Z(_03562_));
 OAI21_X2 _26567_ (.A(_03557_),
    .B1(_03562_),
    .B2(_03097_),
    .ZN(_03563_));
 AOI21_X1 _26568_ (.A(_03178_),
    .B1(_03227_),
    .B2(_03114_),
    .ZN(_03564_));
 OAI222_X2 _26569_ (.A1(_02976_),
    .A2(_03054_),
    .B1(_03093_),
    .B2(_15169_),
    .C1(_03191_),
    .C2(_03122_),
    .ZN(_03565_));
 AOI221_X2 _26570_ (.A(_03166_),
    .B1(_03110_),
    .B2(_03564_),
    .C1(_03565_),
    .C2(_03030_),
    .ZN(_03566_));
 OAI221_X1 _26571_ (.A(_03107_),
    .B1(_03102_),
    .B2(_15172_),
    .C1(_03383_),
    .C2(_02971_),
    .ZN(_03567_));
 NAND3_X1 _26572_ (.A1(_02976_),
    .A2(_03046_),
    .A3(_03047_),
    .ZN(_03568_));
 NAND3_X1 _26573_ (.A1(_02975_),
    .A2(_03116_),
    .A3(_03568_),
    .ZN(_03569_));
 OAI211_X2 _26574_ (.A(_03115_),
    .B(_03173_),
    .C1(_02999_),
    .C2(_03000_),
    .ZN(_03570_));
 NAND3_X1 _26575_ (.A1(_03076_),
    .A2(_03569_),
    .A3(_03570_),
    .ZN(_03571_));
 NAND3_X1 _26576_ (.A1(_03097_),
    .A2(_03567_),
    .A3(_03571_),
    .ZN(_03572_));
 AOI21_X2 _26577_ (.A(_03141_),
    .B1(_03566_),
    .B2(_03572_),
    .ZN(_03573_));
 AOI221_X2 _26578_ (.A(_03540_),
    .B1(_03544_),
    .B2(_03551_),
    .C1(_03573_),
    .C2(_03563_),
    .ZN(_00127_));
 INV_X1 _26579_ (.A(_06340_),
    .ZN(_03574_));
 NOR2_X1 _26580_ (.A1(_03574_),
    .A2(_09730_),
    .ZN(_03575_));
 NOR2_X1 _26581_ (.A1(_06340_),
    .A2(_09728_),
    .ZN(_03576_));
 XNOR2_X2 _26582_ (.A(_08978_),
    .B(_09152_),
    .ZN(_03577_));
 XNOR2_X2 _26583_ (.A(_11856_),
    .B(_03577_),
    .ZN(_03578_));
 XNOR2_X2 _26584_ (.A(_08983_),
    .B(net837),
    .ZN(_03579_));
 XNOR2_X2 _26585_ (.A(_03579_),
    .B(_03578_),
    .ZN(_03580_));
 MUX2_X2 _26586_ (.A(_03575_),
    .B(_03576_),
    .S(_03580_),
    .Z(_03581_));
 OR3_X4 _26587_ (.A1(_06340_),
    .A2(_09856_),
    .A3(_00476_),
    .ZN(_03582_));
 NAND3_X2 _26588_ (.A1(_06340_),
    .A2(_09103_),
    .A3(_00476_),
    .ZN(_03583_));
 NAND2_X4 _26589_ (.A1(_03583_),
    .A2(_03582_),
    .ZN(_03584_));
 NOR2_X4 _26590_ (.A1(_03581_),
    .A2(_03584_),
    .ZN(_03585_));
 INV_X8 _26591_ (.A(net690),
    .ZN(_03586_));
 INV_X4 clone156 (.A(net512),
    .ZN(net156));
 BUF_X16 _26593_ (.A(_03586_),
    .Z(_03588_));
 BUF_X2 rebuffer313 (.A(_03942_),
    .Z(net849));
 XNOR2_X1 _26595_ (.A(\sa00_sr[0] ),
    .B(_03577_),
    .ZN(_03589_));
 NAND3_X1 _26596_ (.A1(_06325_),
    .A2(_09022_),
    .A3(_09019_),
    .ZN(_03590_));
 NOR2_X1 _26597_ (.A1(_06325_),
    .A2(_08971_),
    .ZN(_03591_));
 NAND2_X1 _26598_ (.A1(_09007_),
    .A2(_03591_),
    .ZN(_03592_));
 AOI21_X1 _26599_ (.A(_03589_),
    .B1(_03590_),
    .B2(_03592_),
    .ZN(_03593_));
 XOR2_X1 _26600_ (.A(\sa00_sr[0] ),
    .B(_03577_),
    .Z(_03594_));
 NAND2_X1 _26601_ (.A1(_09019_),
    .A2(_03591_),
    .ZN(_03595_));
 NAND3_X1 _26602_ (.A1(_06325_),
    .A2(_09010_),
    .A3(_09007_),
    .ZN(_03596_));
 AOI21_X1 _26603_ (.A(_03594_),
    .B1(_03595_),
    .B2(_03596_),
    .ZN(_03597_));
 INV_X1 _26604_ (.A(_06325_),
    .ZN(_03598_));
 NAND3_X1 _26605_ (.A1(_03598_),
    .A2(_08972_),
    .A3(_00477_),
    .ZN(_03599_));
 NAND2_X1 _26606_ (.A1(_06325_),
    .A2(_09726_),
    .ZN(_03600_));
 OAI21_X1 _26607_ (.A(_03599_),
    .B1(_03600_),
    .B2(_00477_),
    .ZN(_03601_));
 OR3_X2 _26608_ (.A1(_03593_),
    .A2(_03597_),
    .A3(_03601_),
    .ZN(_03602_));
 BUF_X4 _26609_ (.A(_03602_),
    .Z(_03603_));
 INV_X4 _26610_ (.A(_03603_),
    .ZN(_03604_));
 BUF_X8 _26611_ (.A(_03604_),
    .Z(_03605_));
 BUF_X8 _26612_ (.A(_03605_),
    .Z(_15203_));
 XNOR2_X1 _26613_ (.A(_09088_),
    .B(_09042_),
    .ZN(_03606_));
 INV_X1 _26614_ (.A(net1165),
    .ZN(_03607_));
 NOR3_X1 _26615_ (.A1(_03607_),
    .A2(_11938_),
    .A3(net714),
    .ZN(_03608_));
 NOR3_X1 _26616_ (.A1(net1165),
    .A2(_11841_),
    .A3(net684),
    .ZN(_03609_));
 OAI21_X1 _26617_ (.A(_03606_),
    .B1(_03608_),
    .B2(_03609_),
    .ZN(_03610_));
 XNOR2_X1 _26618_ (.A(_09088_),
    .B(_09044_),
    .ZN(_03611_));
 NOR3_X1 _26619_ (.A1(net1165),
    .A2(_08994_),
    .A3(net714),
    .ZN(_03612_));
 NOR3_X1 _26620_ (.A1(_03607_),
    .A2(_11841_),
    .A3(net684),
    .ZN(_03613_));
 OAI21_X1 _26621_ (.A(_03611_),
    .B1(_03612_),
    .B2(_03613_),
    .ZN(_03614_));
 NAND2_X1 _26622_ (.A1(net1165),
    .A2(_09030_),
    .ZN(_03615_));
 NAND2_X1 _26623_ (.A1(_03607_),
    .A2(_09030_),
    .ZN(_03616_));
 MUX2_X1 _26624_ (.A(_03615_),
    .B(_03616_),
    .S(_00478_),
    .Z(_03617_));
 AND3_X4 _26625_ (.A1(_03610_),
    .A2(_03614_),
    .A3(_03617_),
    .ZN(_03618_));
 INV_X4 _26626_ (.A(_03618_),
    .ZN(_03619_));
 BUF_X4 _26627_ (.A(_03619_),
    .Z(_03620_));
 BUF_X4 _26628_ (.A(_03620_),
    .Z(_03621_));
 BUF_X4 _26629_ (.A(_03621_),
    .Z(_15219_));
 BUF_X4 _26630_ (.A(_03603_),
    .Z(_15194_));
 BUF_X4 _26631_ (.A(_03618_),
    .Z(_03622_));
 BUF_X4 _26632_ (.A(_03622_),
    .Z(_03623_));
 BUF_X4 _26633_ (.A(_03623_),
    .Z(_03624_));
 BUF_X4 _26634_ (.A(_03624_),
    .Z(_15212_));
 OR2_X1 _26635_ (.A1(_09138_),
    .A2(\text_in_r[100] ),
    .ZN(_03625_));
 XNOR2_X2 _26636_ (.A(_09189_),
    .B(_01016_),
    .ZN(_03626_));
 OAI211_X4 _26637_ (.A(_06403_),
    .B(_03625_),
    .C1(_03626_),
    .C2(_09824_),
    .ZN(_03627_));
 INV_X1 _26638_ (.A(_06403_),
    .ZN(_03628_));
 NAND2_X1 _26639_ (.A1(_09824_),
    .A2(\text_in_r[100] ),
    .ZN(_03629_));
 XOR2_X2 _26640_ (.A(_09189_),
    .B(_01016_),
    .Z(_03630_));
 OAI211_X4 _26641_ (.A(_03628_),
    .B(_03629_),
    .C1(_03630_),
    .C2(_09824_),
    .ZN(_03631_));
 NAND2_X4 _26642_ (.A1(_03627_),
    .A2(_03631_),
    .ZN(_03632_));
 CLKBUF_X3 _26643_ (.A(_03632_),
    .Z(_03633_));
 XOR2_X2 _26644_ (.A(_09162_),
    .B(_09165_),
    .Z(_03634_));
 NAND3_X1 _26645_ (.A1(_06417_),
    .A2(_09158_),
    .A3(_03634_),
    .ZN(_03635_));
 NOR2_X1 _26646_ (.A1(_06417_),
    .A2(_09180_),
    .ZN(_03636_));
 NAND2_X1 _26647_ (.A1(_03634_),
    .A2(_03636_),
    .ZN(_03637_));
 MUX2_X2 _26648_ (.A(_03635_),
    .B(_03637_),
    .S(_00996_),
    .Z(_03638_));
 XNOR2_X1 _26649_ (.A(_09162_),
    .B(_09165_),
    .ZN(_03639_));
 NAND2_X1 _26650_ (.A1(_03639_),
    .A2(_03636_),
    .ZN(_03640_));
 NAND3_X1 _26651_ (.A1(_06417_),
    .A2(_09158_),
    .A3(_03639_),
    .ZN(_03641_));
 MUX2_X2 _26652_ (.A(_03640_),
    .B(_03641_),
    .S(_00996_),
    .Z(_03642_));
 OR3_X2 _26653_ (.A1(_06417_),
    .A2(_09803_),
    .A3(\text_in_r[101] ),
    .ZN(_03643_));
 NAND3_X2 _26654_ (.A1(_06417_),
    .A2(_09136_),
    .A3(\text_in_r[101] ),
    .ZN(_03644_));
 AND4_X4 _26655_ (.A1(_03638_),
    .A2(_03642_),
    .A3(_03643_),
    .A4(_03644_),
    .ZN(_03645_));
 BUF_X4 _26656_ (.A(_03645_),
    .Z(_03646_));
 BUF_X4 _26657_ (.A(_03619_),
    .Z(_03647_));
 NOR2_X2 clone2 (.A1(_11851_),
    .A2(net553),
    .ZN(net2));
 INV_X4 _26659_ (.A(_15210_),
    .ZN(_03649_));
 INV_X1 _26660_ (.A(_06386_),
    .ZN(_03650_));
 BUF_X2 _26661_ (.A(\text_in_r[99] ),
    .Z(_03651_));
 NOR2_X1 _26662_ (.A1(_09116_),
    .A2(_03651_),
    .ZN(_03652_));
 XOR2_X2 _26663_ (.A(_09091_),
    .B(_01034_),
    .Z(_03653_));
 AOI211_X4 _26664_ (.A(_03650_),
    .B(_03652_),
    .C1(_03653_),
    .C2(_09175_),
    .ZN(_03654_));
 BUF_X8 _26665_ (.A(_03654_),
    .Z(_03655_));
 INV_X1 _26666_ (.A(_03651_),
    .ZN(_03656_));
 NOR2_X1 _26667_ (.A1(net594),
    .A2(_03656_),
    .ZN(_03657_));
 XNOR2_X2 _26668_ (.A(_09091_),
    .B(_01034_),
    .ZN(_03658_));
 AOI211_X4 _26669_ (.A(_06386_),
    .B(_03657_),
    .C1(_03658_),
    .C2(_11191_),
    .ZN(_03659_));
 BUF_X8 _26670_ (.A(_03659_),
    .Z(_03660_));
 NOR3_X4 _26671_ (.A1(_03649_),
    .A2(_03655_),
    .A3(_03660_),
    .ZN(_03661_));
 NAND2_X1 _26672_ (.A1(_08996_),
    .A2(_03656_),
    .ZN(_03662_));
 OAI211_X4 _26673_ (.A(_06386_),
    .B(_03662_),
    .C1(_03658_),
    .C2(_09824_),
    .ZN(_03663_));
 BUF_X8 _26674_ (.A(_03663_),
    .Z(_03664_));
 NAND2_X1 _26675_ (.A1(_09135_),
    .A2(_03651_),
    .ZN(_03665_));
 OAI211_X4 _26676_ (.A(_03650_),
    .B(_03665_),
    .C1(_03653_),
    .C2(_09824_),
    .ZN(_03666_));
 BUF_X8 _26677_ (.A(_03666_),
    .Z(_03667_));
 AOI211_X2 _26678_ (.A(net560),
    .B(_03584_),
    .C1(_03664_),
    .C2(_03667_),
    .ZN(_03668_));
 OAI21_X4 _26679_ (.A(_03647_),
    .B1(_03668_),
    .B2(_03661_),
    .ZN(_03669_));
 NAND3_X2 _26680_ (.A1(_03622_),
    .A2(_03664_),
    .A3(_03667_),
    .ZN(_03670_));
 BUF_X4 _26681_ (.A(_03670_),
    .Z(_03671_));
 BUF_X4 _26682_ (.A(_15197_),
    .Z(_03672_));
 INV_X4 _26683_ (.A(_03672_),
    .ZN(_03673_));
 BUF_X8 _26684_ (.A(_03673_),
    .Z(_03674_));
 NOR2_X4 _26685_ (.A1(_03654_),
    .A2(_03659_),
    .ZN(_03675_));
 BUF_X4 _26686_ (.A(_03675_),
    .Z(_03676_));
 BUF_X4 _26687_ (.A(_03676_),
    .Z(_03677_));
 OAI221_X2 _26688_ (.A(_03669_),
    .B1(_03671_),
    .B2(net155),
    .C1(_15194_),
    .C2(_03677_),
    .ZN(_03678_));
 NAND2_X1 _26689_ (.A1(_06340_),
    .A2(_11192_),
    .ZN(_03679_));
 NAND2_X1 _26690_ (.A1(_03574_),
    .A2(_11192_),
    .ZN(_03680_));
 MUX2_X2 _26691_ (.A(_03679_),
    .B(_03680_),
    .S(net747),
    .Z(_03681_));
 AND2_X2 _26692_ (.A1(_03582_),
    .A2(_03583_),
    .ZN(_03682_));
 OAI211_X4 _26693_ (.A(_03681_),
    .B(_03682_),
    .C1(_03655_),
    .C2(_03660_),
    .ZN(_03683_));
 NOR2_X2 _26694_ (.A1(_03605_),
    .A2(_03618_),
    .ZN(_03684_));
 AOI21_X1 _26695_ (.A(_03646_),
    .B1(_03683_),
    .B2(_03684_),
    .ZN(_03685_));
 BUF_X4 _26696_ (.A(_03623_),
    .Z(_03686_));
 BUF_X4 _26697_ (.A(_03686_),
    .Z(_03687_));
 BUF_X4 _26698_ (.A(_03664_),
    .Z(_03688_));
 BUF_X4 _26699_ (.A(_03667_),
    .Z(_03689_));
 NAND3_X1 _26700_ (.A1(net744),
    .A2(_03688_),
    .A3(_03689_),
    .ZN(_03690_));
 OAI22_X4 _26701_ (.A1(net560),
    .A2(_03584_),
    .B1(_03654_),
    .B2(_03659_),
    .ZN(_03691_));
 NAND3_X1 _26702_ (.A1(_03687_),
    .A2(_03690_),
    .A3(_03691_),
    .ZN(_03692_));
 AOI221_X2 _26703_ (.A(_03633_),
    .B1(_03678_),
    .B2(_03646_),
    .C1(_03685_),
    .C2(_03692_),
    .ZN(_03693_));
 XNOR2_X2 _26704_ (.A(_09014_),
    .B(_11897_),
    .ZN(_03694_));
 XNOR2_X2 _26705_ (.A(_09151_),
    .B(_03694_),
    .ZN(_03695_));
 MUX2_X2 _26706_ (.A(\text_in_r[103] ),
    .B(_03695_),
    .S(_11192_),
    .Z(_03696_));
 XNOR2_X2 _26707_ (.A(_06439_),
    .B(_03696_),
    .ZN(_03697_));
 CLKBUF_X3 _26708_ (.A(_03697_),
    .Z(_03698_));
 BUF_X8 clone154 (.A(_03716_),
    .Z(net154));
 INV_X8 _26710_ (.A(net847),
    .ZN(_03700_));
 NOR3_X4 _26711_ (.A1(_03620_),
    .A2(_03655_),
    .A3(_03660_),
    .ZN(_03701_));
 NAND4_X4 _26712_ (.A1(_03681_),
    .A2(_03682_),
    .A3(_03663_),
    .A4(_03666_),
    .ZN(_03702_));
 AOI22_X1 _26713_ (.A1(_03700_),
    .A2(_03701_),
    .B1(_03702_),
    .B2(_03684_),
    .ZN(_03703_));
 NAND2_X2 _26714_ (.A1(_03632_),
    .A2(_03645_),
    .ZN(_03704_));
 BUF_X4 _26715_ (.A(_03704_),
    .Z(_03705_));
 AND2_X1 _26716_ (.A1(_03627_),
    .A2(_03631_),
    .ZN(_03706_));
 CLKBUF_X3 _26717_ (.A(_03706_),
    .Z(_03707_));
 BUF_X4 _26718_ (.A(_03707_),
    .Z(_03708_));
 NAND2_X4 _26719_ (.A1(_03663_),
    .A2(_03666_),
    .ZN(_03709_));
 NOR2_X4 _26720_ (.A1(_03603_),
    .A2(_03619_),
    .ZN(_03710_));
 AOI211_X2 _26721_ (.A(_03709_),
    .B(_03684_),
    .C1(_03710_),
    .C2(_03586_),
    .ZN(_03711_));
 OR2_X1 _26722_ (.A1(_03708_),
    .A2(_03711_),
    .ZN(_03712_));
 NAND4_X4 _26723_ (.A1(_03638_),
    .A2(_03642_),
    .A3(_03643_),
    .A4(_03644_),
    .ZN(_03713_));
 BUF_X4 _26724_ (.A(_03713_),
    .Z(_03714_));
 BUF_X4 _26725_ (.A(_03714_),
    .Z(_03715_));
 BUF_X8 _26726_ (.A(_03585_),
    .Z(_03716_));
 NOR2_X1 _26727_ (.A1(net153),
    .A2(_03686_),
    .ZN(_03717_));
 BUF_X4 _26728_ (.A(_03709_),
    .Z(_03718_));
 CLKBUF_X3 _26729_ (.A(_03718_),
    .Z(_03719_));
 BUF_X4 _26730_ (.A(_03621_),
    .Z(_03720_));
 BUF_X2 _26731_ (.A(_15198_),
    .Z(_03721_));
 BUF_X4 _26732_ (.A(_03721_),
    .Z(_03722_));
 OAI21_X1 _26733_ (.A(_03719_),
    .B1(_03720_),
    .B2(_03722_),
    .ZN(_03723_));
 OAI21_X1 _26734_ (.A(_03715_),
    .B1(_03717_),
    .B2(_03723_),
    .ZN(_03724_));
 OAI221_X1 _26735_ (.A(_03698_),
    .B1(_03703_),
    .B2(_03705_),
    .C1(_03712_),
    .C2(_03724_),
    .ZN(_03725_));
 TAPCELL_X1 PHY_EDGE_ROW_1_Right_1 ();
 BUF_X4 _26737_ (.A(_03709_),
    .Z(_03727_));
 NAND2_X1 _26738_ (.A1(net943),
    .A2(_03727_),
    .ZN(_03728_));
 OAI221_X1 _26739_ (.A(_03708_),
    .B1(_03671_),
    .B2(net155),
    .C1(_03728_),
    .C2(_03621_),
    .ZN(_03729_));
 NOR3_X4 _26740_ (.A1(_03605_),
    .A2(_03654_),
    .A3(_03659_),
    .ZN(_03730_));
 NAND2_X1 _26741_ (.A1(_03632_),
    .A2(_03730_),
    .ZN(_03731_));
 BUF_X4 _26742_ (.A(_15201_),
    .Z(_03732_));
 NOR2_X1 _26743_ (.A1(_03732_),
    .A2(_03677_),
    .ZN(_03733_));
 NOR2_X1 _26744_ (.A1(_03687_),
    .A2(_03733_),
    .ZN(_03734_));
 AOI221_X1 _26745_ (.A(_03646_),
    .B1(_03712_),
    .B2(_03729_),
    .C1(_03731_),
    .C2(_03734_),
    .ZN(_03735_));
 XOR2_X2 _26746_ (.A(_06439_),
    .B(_03696_),
    .Z(_03736_));
 CLKBUF_X3 _26747_ (.A(_03727_),
    .Z(_03737_));
 BUF_X8 _26748_ (.A(_03672_),
    .Z(_03738_));
 NAND2_X1 _26749_ (.A1(_03738_),
    .A2(_03647_),
    .ZN(_03739_));
 OAI21_X4 _26750_ (.A(_03622_),
    .B1(_03584_),
    .B2(_03581_),
    .ZN(_03740_));
 NAND3_X1 _26751_ (.A1(_03737_),
    .A2(_03739_),
    .A3(_03740_),
    .ZN(_03741_));
 BUF_X4 _26752_ (.A(_03677_),
    .Z(_03742_));
 BUF_X4 _26753_ (.A(_15204_),
    .Z(_03743_));
 NOR2_X1 _26754_ (.A1(_03743_),
    .A2(_03686_),
    .ZN(_03744_));
 OAI21_X1 _26755_ (.A(_03742_),
    .B1(_03710_),
    .B2(_03744_),
    .ZN(_03745_));
 NAND2_X1 _26756_ (.A1(_03741_),
    .A2(_03745_),
    .ZN(_03746_));
 NAND2_X4 _26757_ (.A1(_03708_),
    .A2(_03645_),
    .ZN(_03747_));
 OAI21_X4 _26758_ (.A(_03622_),
    .B1(_03655_),
    .B2(_03660_),
    .ZN(_03748_));
 OAI22_X1 _26759_ (.A1(_03732_),
    .A2(_03671_),
    .B1(_03748_),
    .B2(_03722_),
    .ZN(_03749_));
 AOI21_X4 _26760_ (.A(_03622_),
    .B1(_03688_),
    .B2(_03689_),
    .ZN(_03750_));
 BUF_X4 clone157 (.A(_03586_),
    .Z(net157));
 AOI21_X1 _26762_ (.A(_03749_),
    .B1(_03750_),
    .B2(net746),
    .ZN(_03752_));
 OAI221_X1 _26763_ (.A(_03736_),
    .B1(_03705_),
    .B2(_03746_),
    .C1(_03747_),
    .C2(_03752_),
    .ZN(_03753_));
 OAI22_X1 _26764_ (.A1(_03725_),
    .A2(_03693_),
    .B1(_03735_),
    .B2(_03753_),
    .ZN(_03754_));
 AOI21_X4 _26765_ (.A(_03721_),
    .B1(_03664_),
    .B2(_03667_),
    .ZN(_03755_));
 AOI21_X1 _26766_ (.A(_03755_),
    .B1(_03730_),
    .B2(net156),
    .ZN(_03756_));
 NOR3_X2 _26767_ (.A1(_03622_),
    .A2(_03655_),
    .A3(_03660_),
    .ZN(_03757_));
 BUF_X4 _26768_ (.A(_03757_),
    .Z(_03758_));
 AOI221_X2 _26769_ (.A(_03705_),
    .B1(_03756_),
    .B2(_03687_),
    .C1(_03758_),
    .C2(net944),
    .ZN(_03759_));
 CLKBUF_X3 _26770_ (.A(_03736_),
    .Z(_03760_));
 CLKBUF_X3 _26771_ (.A(_03715_),
    .Z(_03761_));
 BUF_X4 _26772_ (.A(_03707_),
    .Z(_03762_));
 BUF_X4 _26773_ (.A(_03762_),
    .Z(_03763_));
 OAI21_X2 _26774_ (.A(_03603_),
    .B1(_03584_),
    .B2(_03581_),
    .ZN(_03764_));
 OAI21_X2 _26775_ (.A(_03718_),
    .B1(_03764_),
    .B2(_03647_),
    .ZN(_03765_));
 INV_X2 _26776_ (.A(_03743_),
    .ZN(_03766_));
 NOR2_X1 _26777_ (.A1(_03766_),
    .A2(_03623_),
    .ZN(_03767_));
 NAND3_X2 _26778_ (.A1(_03722_),
    .A2(_03688_),
    .A3(_03689_),
    .ZN(_03768_));
 OAI221_X2 _26779_ (.A(_03763_),
    .B1(_03765_),
    .B2(_03767_),
    .C1(_03768_),
    .C2(_15219_),
    .ZN(_03769_));
 OAI21_X1 _26780_ (.A(_03760_),
    .B1(_03761_),
    .B2(_03769_),
    .ZN(_03770_));
 BUF_X4 _26781_ (.A(_03646_),
    .Z(_03771_));
 BUF_X4 _26782_ (.A(_03632_),
    .Z(_03772_));
 INV_X2 _26783_ (.A(net745),
    .ZN(_03773_));
 OAI221_X1 _26784_ (.A(_03772_),
    .B1(_03748_),
    .B2(_03764_),
    .C1(_03671_),
    .C2(_03773_),
    .ZN(_03774_));
 OR2_X1 _26785_ (.A1(_03730_),
    .A2(_03755_),
    .ZN(_03775_));
 AOI21_X1 _26786_ (.A(_03774_),
    .B1(_03775_),
    .B2(_03720_),
    .ZN(_03776_));
 OAI21_X4 _26787_ (.A(net693),
    .B1(_03655_),
    .B2(_03660_),
    .ZN(_03777_));
 NAND2_X2 _26788_ (.A1(_03620_),
    .A2(_03707_),
    .ZN(_03778_));
 NAND2_X1 _26789_ (.A1(_03707_),
    .A2(_03676_),
    .ZN(_03779_));
 INV_X1 _26790_ (.A(_15217_),
    .ZN(_03780_));
 OAI22_X1 _26791_ (.A1(_03777_),
    .A2(_03778_),
    .B1(_03779_),
    .B2(_03780_),
    .ZN(_03781_));
 NOR3_X1 _26792_ (.A1(_03700_),
    .A2(_03762_),
    .A3(_03765_),
    .ZN(_03782_));
 NOR4_X2 _26793_ (.A1(_03771_),
    .A2(_03776_),
    .A3(_03781_),
    .A4(_03782_),
    .ZN(_03783_));
 OAI211_X4 _26794_ (.A(_03627_),
    .B(_03631_),
    .C1(_03655_),
    .C2(_03660_),
    .ZN(_03784_));
 NAND3_X1 _26795_ (.A1(_03738_),
    .A2(_03687_),
    .A3(_03715_),
    .ZN(_03785_));
 NAND2_X2 _26796_ (.A1(_03605_),
    .A2(_03647_),
    .ZN(_03786_));
 BUF_X16 _26797_ (.A(_03716_),
    .Z(_15195_));
 BUF_X4 _26798_ (.A(_03647_),
    .Z(_03787_));
 AOI21_X1 _26799_ (.A(_03787_),
    .B1(_03646_),
    .B2(_15194_),
    .ZN(_03788_));
 OAI221_X1 _26800_ (.A(_03785_),
    .B1(_03786_),
    .B2(_03715_),
    .C1(net154),
    .C2(_03788_),
    .ZN(_03789_));
 NOR2_X1 _26801_ (.A1(_03784_),
    .A2(_03789_),
    .ZN(_03790_));
 NAND2_X1 _26802_ (.A1(_03766_),
    .A2(_03742_),
    .ZN(_03791_));
 AOI21_X4 _26803_ (.A(_03674_),
    .B1(_03688_),
    .B2(_03689_),
    .ZN(_03792_));
 NOR2_X4 _26804_ (.A1(_03792_),
    .A2(_03621_),
    .ZN(_03793_));
 BUF_X4 _26805_ (.A(_03654_),
    .Z(_03794_));
 BUF_X4 _26806_ (.A(_03659_),
    .Z(_03795_));
 NOR3_X2 _26807_ (.A1(net745),
    .A2(_03794_),
    .A3(_03795_),
    .ZN(_03796_));
 OAI21_X4 _26808_ (.A(_03604_),
    .B1(_03584_),
    .B2(net561),
    .ZN(_03797_));
 AOI21_X1 _26809_ (.A(_03796_),
    .B1(_03797_),
    .B2(_03737_),
    .ZN(_03798_));
 AOI22_X4 _26810_ (.A1(_03793_),
    .A2(_03791_),
    .B1(_03798_),
    .B2(_03720_),
    .ZN(_03799_));
 NOR2_X2 _26811_ (.A1(_03705_),
    .A2(_03799_),
    .ZN(_03800_));
 NOR2_X2 _26812_ (.A1(_03674_),
    .A2(_03670_),
    .ZN(_03801_));
 OAI21_X4 _26813_ (.A(_03620_),
    .B1(_03655_),
    .B2(_03660_),
    .ZN(_03802_));
 NOR2_X1 _26814_ (.A1(_03743_),
    .A2(_03802_),
    .ZN(_03803_));
 NAND2_X4 _26815_ (.A1(_03632_),
    .A2(_03713_),
    .ZN(_03804_));
 NAND3_X4 _26816_ (.A1(_03619_),
    .A2(_03664_),
    .A3(_03667_),
    .ZN(_03805_));
 AOI21_X1 _26817_ (.A(net745),
    .B1(_03748_),
    .B2(_03805_),
    .ZN(_03806_));
 OR4_X1 _26818_ (.A1(_03801_),
    .A2(_03803_),
    .A3(_03804_),
    .A4(_03806_),
    .ZN(_03807_));
 NOR2_X2 _26819_ (.A1(_03772_),
    .A2(_03718_),
    .ZN(_03808_));
 AOI21_X1 _26820_ (.A(_03710_),
    .B1(_15194_),
    .B2(_15195_),
    .ZN(_03809_));
 NAND2_X1 _26821_ (.A1(_03787_),
    .A2(_03715_),
    .ZN(_03810_));
 OAI221_X2 _26822_ (.A(_03808_),
    .B1(_03809_),
    .B2(_03715_),
    .C1(_03810_),
    .C2(_03738_),
    .ZN(_03811_));
 NAND3_X1 _26823_ (.A1(_03698_),
    .A2(_03807_),
    .A3(_03811_),
    .ZN(_03812_));
 OAI33_X1 _26824_ (.A1(_03759_),
    .A2(_03770_),
    .A3(_03783_),
    .B1(_03800_),
    .B2(_03790_),
    .B3(_03812_),
    .ZN(_03813_));
 XNOR2_X1 _26825_ (.A(_09166_),
    .B(_09154_),
    .ZN(_03814_));
 XNOR2_X2 _26826_ (.A(_09069_),
    .B(_03814_),
    .ZN(_03815_));
 MUX2_X2 _26827_ (.A(\text_in_r[102] ),
    .B(_03815_),
    .S(_11207_),
    .Z(_03816_));
 XNOR2_X2 _26828_ (.A(_06431_),
    .B(_03816_),
    .ZN(_03817_));
 BUF_X4 _26829_ (.A(_03817_),
    .Z(_03818_));
 BUF_X4 _26830_ (.A(_03818_),
    .Z(_03819_));
 MUX2_X1 _26831_ (.A(_03754_),
    .B(_03813_),
    .S(_03819_),
    .Z(_00128_));
 CLKBUF_X3 _26832_ (.A(_03771_),
    .Z(_03820_));
 XOR2_X2 _26833_ (.A(_06431_),
    .B(_03816_),
    .Z(_03821_));
 NAND2_X2 _26834_ (.A1(_03708_),
    .A2(_03714_),
    .ZN(_03822_));
 NAND3_X2 _26835_ (.A1(_03738_),
    .A2(_03688_),
    .A3(_03689_),
    .ZN(_03823_));
 OAI21_X2 _26836_ (.A(net745),
    .B1(_03655_),
    .B2(_03660_),
    .ZN(_03824_));
 NAND3_X1 _26837_ (.A1(_03624_),
    .A2(_03823_),
    .A3(_03824_),
    .ZN(_03825_));
 AOI21_X4 _26838_ (.A(_03603_),
    .B1(_03664_),
    .B2(_03667_),
    .ZN(_03826_));
 NOR3_X4 _26839_ (.A1(_03700_),
    .A2(_03654_),
    .A3(_03659_),
    .ZN(_03827_));
 OAI21_X1 _26840_ (.A(_03787_),
    .B1(_03826_),
    .B2(_03827_),
    .ZN(_03828_));
 AND2_X1 _26841_ (.A1(_03825_),
    .A2(_03828_),
    .ZN(_03829_));
 NOR2_X4 _26842_ (.A1(_03605_),
    .A2(_03619_),
    .ZN(_03830_));
 OAI21_X1 _26843_ (.A(_03748_),
    .B1(_03718_),
    .B2(_03716_),
    .ZN(_03831_));
 AOI222_X2 _26844_ (.A1(net155),
    .A2(_03750_),
    .B1(_03830_),
    .B2(_03742_),
    .C1(_03831_),
    .C2(_15203_),
    .ZN(_03832_));
 OAI221_X2 _26845_ (.A(_03821_),
    .B1(_03822_),
    .B2(_03829_),
    .C1(_03832_),
    .C2(_03804_),
    .ZN(_03833_));
 MUX2_X1 _26846_ (.A(_03674_),
    .B(_03649_),
    .S(_03623_),
    .Z(_03834_));
 OAI21_X2 _26847_ (.A(_03772_),
    .B1(_03834_),
    .B2(_03737_),
    .ZN(_03835_));
 AOI221_X2 _26848_ (.A(_03676_),
    .B1(_03830_),
    .B2(_03586_),
    .C1(_03647_),
    .C2(_03700_),
    .ZN(_03836_));
 OAI21_X1 _26849_ (.A(_03715_),
    .B1(_03836_),
    .B2(_03835_),
    .ZN(_03837_));
 NAND2_X1 _26850_ (.A1(_03700_),
    .A2(_03750_),
    .ZN(_03838_));
 AOI21_X4 _26851_ (.A(_03620_),
    .B1(_03688_),
    .B2(_03689_),
    .ZN(_03839_));
 OAI21_X1 _26852_ (.A(net850),
    .B1(_03839_),
    .B2(_03758_),
    .ZN(_03840_));
 AOI21_X1 _26853_ (.A(_03633_),
    .B1(_03838_),
    .B2(_03840_),
    .ZN(_03841_));
 OAI21_X1 _26854_ (.A(_03819_),
    .B1(_03837_),
    .B2(_03841_),
    .ZN(_03842_));
 AOI21_X1 _26855_ (.A(_03820_),
    .B1(_03833_),
    .B2(_03842_),
    .ZN(_03843_));
 OR2_X1 _26856_ (.A1(_03837_),
    .A2(_03841_),
    .ZN(_03844_));
 CLKBUF_X3 _26857_ (.A(_03686_),
    .Z(_03845_));
 NAND3_X2 _26858_ (.A1(_03605_),
    .A2(_03688_),
    .A3(_03689_),
    .ZN(_03846_));
 AOI21_X4 _26859_ (.A(_03605_),
    .B1(_03664_),
    .B2(_03667_),
    .ZN(_03847_));
 OAI21_X1 _26860_ (.A(_03847_),
    .B1(_03762_),
    .B2(net850),
    .ZN(_03848_));
 AOI21_X1 _26861_ (.A(_03845_),
    .B1(_03846_),
    .B2(_03848_),
    .ZN(_03849_));
 OAI21_X2 _26862_ (.A(_03732_),
    .B1(_03794_),
    .B2(_03795_),
    .ZN(_03850_));
 AOI21_X1 _26863_ (.A(_03633_),
    .B1(_03823_),
    .B2(_03850_),
    .ZN(_03851_));
 AOI21_X1 _26864_ (.A(_03849_),
    .B1(_03851_),
    .B2(_15212_),
    .ZN(_03852_));
 CLKBUF_X3 _26865_ (.A(_03772_),
    .Z(_03853_));
 NOR2_X1 _26866_ (.A1(_03603_),
    .A2(_03623_),
    .ZN(_03854_));
 OAI21_X2 _26867_ (.A(_03605_),
    .B1(_03794_),
    .B2(_03795_),
    .ZN(_03855_));
 AOI21_X1 _26868_ (.A(net157),
    .B1(_03855_),
    .B2(_03805_),
    .ZN(_03856_));
 OAI21_X1 _26869_ (.A(_03853_),
    .B1(_03854_),
    .B2(_03856_),
    .ZN(_03857_));
 AND4_X1 _26870_ (.A1(_03819_),
    .A2(_03844_),
    .A3(_03852_),
    .A4(_03857_),
    .ZN(_03858_));
 AOI21_X1 _26871_ (.A(_03633_),
    .B1(_03826_),
    .B2(_03588_),
    .ZN(_03859_));
 OAI221_X1 _26872_ (.A(_03859_),
    .B1(_03661_),
    .B2(_03845_),
    .C1(net195),
    .C2(_03671_),
    .ZN(_03860_));
 NAND3_X4 _26873_ (.A1(_03673_),
    .A2(_03664_),
    .A3(_03667_),
    .ZN(_03861_));
 AOI21_X1 _26874_ (.A(_03720_),
    .B1(_03861_),
    .B2(_03850_),
    .ZN(_03862_));
 AOI21_X1 _26875_ (.A(_03862_),
    .B1(_03758_),
    .B2(_03797_),
    .ZN(_03863_));
 BUF_X4 _26876_ (.A(_03708_),
    .Z(_03864_));
 BUF_X4 _26877_ (.A(_03864_),
    .Z(_03865_));
 OAI21_X1 _26878_ (.A(_03860_),
    .B1(_03863_),
    .B2(_03865_),
    .ZN(_03866_));
 OAI21_X1 _26879_ (.A(_03760_),
    .B1(_03833_),
    .B2(_03866_),
    .ZN(_03867_));
 OR2_X4 _26880_ (.A1(_03827_),
    .A2(_03619_),
    .ZN(_03868_));
 AND2_X1 _26881_ (.A1(_03691_),
    .A2(_03702_),
    .ZN(_03869_));
 OAI221_X1 _26882_ (.A(_03761_),
    .B1(_03847_),
    .B2(_03868_),
    .C1(_03869_),
    .C2(_15212_),
    .ZN(_03870_));
 NAND2_X1 _26883_ (.A1(net156),
    .A2(_03676_),
    .ZN(_03871_));
 OR2_X1 _26884_ (.A1(_03830_),
    .A2(_03854_),
    .ZN(_03872_));
 AOI21_X1 _26885_ (.A(_03830_),
    .B1(_15219_),
    .B2(net745),
    .ZN(_03873_));
 OAI221_X1 _26886_ (.A(_03771_),
    .B1(_03871_),
    .B2(_03872_),
    .C1(_03873_),
    .C2(_03742_),
    .ZN(_03874_));
 NAND3_X1 _26887_ (.A1(_03865_),
    .A2(_03870_),
    .A3(_03874_),
    .ZN(_03875_));
 AOI221_X2 _26888_ (.A(_03675_),
    .B1(_03710_),
    .B2(_03586_),
    .C1(_03620_),
    .C2(net187),
    .ZN(_03876_));
 NOR2_X2 _26889_ (.A1(_03762_),
    .A2(_03876_),
    .ZN(_03877_));
 NAND2_X1 _26890_ (.A1(_03714_),
    .A2(_03677_),
    .ZN(_03878_));
 OAI21_X1 _26891_ (.A(_03877_),
    .B1(_03878_),
    .B2(_15220_),
    .ZN(_03879_));
 AOI21_X1 _26892_ (.A(_03821_),
    .B1(_03875_),
    .B2(_03879_),
    .ZN(_03880_));
 OAI21_X1 _26893_ (.A(_03861_),
    .B1(_03855_),
    .B2(_03716_),
    .ZN(_03881_));
 AOI221_X2 _26894_ (.A(_03804_),
    .B1(_03881_),
    .B2(_03686_),
    .C1(_03750_),
    .C2(_15194_),
    .ZN(_03882_));
 OAI21_X2 _26895_ (.A(net744),
    .B1(_03794_),
    .B2(_03795_),
    .ZN(_03883_));
 NOR3_X4 _26896_ (.A1(net693),
    .A2(_03654_),
    .A3(_03659_),
    .ZN(_03884_));
 NOR2_X4 _26897_ (.A1(_03647_),
    .A2(_03884_),
    .ZN(_03885_));
 OR2_X1 _26898_ (.A1(_03721_),
    .A2(_03675_),
    .ZN(_03886_));
 OAI21_X2 _26899_ (.A(_03886_),
    .B1(_03797_),
    .B2(_03727_),
    .ZN(_03887_));
 AOI221_X2 _26900_ (.A(_03822_),
    .B1(_03883_),
    .B2(_03885_),
    .C1(_03887_),
    .C2(_03787_),
    .ZN(_03888_));
 NOR3_X4 _26901_ (.A1(_03732_),
    .A2(_03794_),
    .A3(_03795_),
    .ZN(_03889_));
 OAI21_X1 _26902_ (.A(_03624_),
    .B1(_03826_),
    .B2(_03889_),
    .ZN(_03890_));
 NOR2_X2 _26903_ (.A1(net745),
    .A2(_03675_),
    .ZN(_03891_));
 OAI21_X1 _26904_ (.A(_03621_),
    .B1(_03718_),
    .B2(net154),
    .ZN(_03892_));
 OAI21_X1 _26905_ (.A(_03890_),
    .B1(_03891_),
    .B2(_03892_),
    .ZN(_03893_));
 BUF_X4 _26906_ (.A(_03676_),
    .Z(_03894_));
 AOI21_X1 _26907_ (.A(_03755_),
    .B1(_03894_),
    .B2(net745),
    .ZN(_03895_));
 NOR2_X1 _26908_ (.A1(_03686_),
    .A2(_03884_),
    .ZN(_03896_));
 OAI21_X2 _26909_ (.A(_03603_),
    .B1(_03655_),
    .B2(_03660_),
    .ZN(_03897_));
 AOI22_X1 _26910_ (.A1(_03687_),
    .A2(_03895_),
    .B1(_03896_),
    .B2(_03897_),
    .ZN(_03898_));
 OAI22_X1 _26911_ (.A1(_03705_),
    .A2(_03893_),
    .B1(_03898_),
    .B2(_03747_),
    .ZN(_03899_));
 NOR4_X1 _26912_ (.A1(_03899_),
    .A2(_03882_),
    .A3(_03888_),
    .A4(_03819_),
    .ZN(_03900_));
 OAI33_X1 _26913_ (.A1(_03858_),
    .A2(_03843_),
    .A3(_03867_),
    .B1(_03880_),
    .B2(_03900_),
    .B3(_03760_),
    .ZN(_00129_));
 NAND3_X1 _26914_ (.A1(net195),
    .A2(_15219_),
    .A3(_03855_),
    .ZN(_03901_));
 OAI221_X1 _26915_ (.A(_03853_),
    .B1(_03730_),
    .B2(_03901_),
    .C1(_03671_),
    .C2(net152),
    .ZN(_03902_));
 AOI21_X4 _26916_ (.A(_03621_),
    .B1(net1036),
    .B2(_03846_),
    .ZN(_03903_));
 AOI21_X1 _26917_ (.A(_15212_),
    .B1(_03683_),
    .B2(_03768_),
    .ZN(_03904_));
 OAI21_X1 _26918_ (.A(_03865_),
    .B1(_03903_),
    .B2(_03904_),
    .ZN(_03905_));
 NAND3_X1 _26919_ (.A1(_03820_),
    .A2(_03902_),
    .A3(_03905_),
    .ZN(_03906_));
 MUX2_X1 _26920_ (.A(_03649_),
    .B(_03700_),
    .S(_03618_),
    .Z(_03907_));
 OAI21_X2 _26921_ (.A(_03714_),
    .B1(_03907_),
    .B2(_03784_),
    .ZN(_03908_));
 NAND2_X1 _26922_ (.A1(net195),
    .A2(_03786_),
    .ZN(_03909_));
 AOI21_X1 _26923_ (.A(_03908_),
    .B1(_03909_),
    .B2(_03808_),
    .ZN(_03910_));
 NAND2_X1 _26924_ (.A1(_03853_),
    .A2(_03741_),
    .ZN(_03911_));
 NAND2_X2 _26925_ (.A1(net156),
    .A2(_03830_),
    .ZN(_03912_));
 BUF_X4 _26926_ (.A(_03622_),
    .Z(_03913_));
 NOR2_X1 _26927_ (.A1(_03732_),
    .A2(_03913_),
    .ZN(_03914_));
 INV_X1 _26928_ (.A(_03914_),
    .ZN(_03915_));
 AOI21_X2 _26929_ (.A(_03737_),
    .B1(_03912_),
    .B2(_03915_),
    .ZN(_03916_));
 OAI21_X1 _26930_ (.A(_03910_),
    .B1(_03911_),
    .B2(_03916_),
    .ZN(_03917_));
 NOR2_X1 _26931_ (.A1(_03760_),
    .A2(_03821_),
    .ZN(_03918_));
 NAND3_X1 _26932_ (.A1(_03906_),
    .A2(_03917_),
    .A3(_03918_),
    .ZN(_03919_));
 INV_X1 _26933_ (.A(_15220_),
    .ZN(_03920_));
 AOI21_X1 _26934_ (.A(_03762_),
    .B1(_03737_),
    .B2(_03920_),
    .ZN(_03921_));
 OAI21_X1 _26935_ (.A(_03740_),
    .B1(_15203_),
    .B2(net850),
    .ZN(_03922_));
 OAI21_X1 _26936_ (.A(_03921_),
    .B1(_03922_),
    .B2(_03719_),
    .ZN(_03923_));
 NAND2_X1 _26937_ (.A1(_03623_),
    .A2(_03707_),
    .ZN(_03924_));
 OAI21_X1 _26938_ (.A(_03691_),
    .B1(_03727_),
    .B2(_03743_),
    .ZN(_03925_));
 NOR2_X1 _26939_ (.A1(_03924_),
    .A2(_03925_),
    .ZN(_03926_));
 AOI21_X1 _26940_ (.A(_03778_),
    .B1(_03861_),
    .B2(_03824_),
    .ZN(_03927_));
 NOR3_X1 _26941_ (.A1(_03646_),
    .A2(_03926_),
    .A3(_03927_),
    .ZN(_03928_));
 NOR2_X1 _26942_ (.A1(net693),
    .A2(_03618_),
    .ZN(_03929_));
 NOR2_X1 _26943_ (.A1(_03709_),
    .A2(_03929_),
    .ZN(_03930_));
 AOI221_X1 _26944_ (.A(_03708_),
    .B1(_03912_),
    .B2(_03930_),
    .C1(_03727_),
    .C2(_15217_),
    .ZN(_03931_));
 AOI22_X2 _26945_ (.A1(_03681_),
    .A2(_03682_),
    .B1(_03688_),
    .B2(_03689_),
    .ZN(_03932_));
 NOR3_X1 _26946_ (.A1(net560),
    .A2(_03584_),
    .A3(_03622_),
    .ZN(_03933_));
 OAI21_X1 _26947_ (.A(_03738_),
    .B1(_03932_),
    .B2(_03933_),
    .ZN(_03934_));
 NOR3_X4 _26948_ (.A1(_03603_),
    .A2(_03794_),
    .A3(_03795_),
    .ZN(_03935_));
 OAI221_X1 _26949_ (.A(_03934_),
    .B1(_03935_),
    .B2(_03740_),
    .C1(_03702_),
    .C2(_03710_),
    .ZN(_03936_));
 AOI21_X1 _26950_ (.A(_03931_),
    .B1(_03936_),
    .B2(_03763_),
    .ZN(_03937_));
 AOI221_X2 _26951_ (.A(_03818_),
    .B1(_03923_),
    .B2(_03928_),
    .C1(_03937_),
    .C2(_03771_),
    .ZN(_03938_));
 NOR3_X1 _26952_ (.A1(_06386_),
    .A2(_03658_),
    .A3(_03657_),
    .ZN(_03939_));
 NOR2_X1 _26953_ (.A1(_03650_),
    .A2(_09136_),
    .ZN(_03940_));
 AOI21_X2 _26954_ (.A(_03939_),
    .B1(_03940_),
    .B2(_03658_),
    .ZN(_03941_));
 OR2_X4 _26955_ (.A1(_03721_),
    .A2(_15201_),
    .ZN(_03942_));
 NOR3_X1 _26956_ (.A1(_06386_),
    .A2(_09158_),
    .A3(_03651_),
    .ZN(_03943_));
 AOI21_X2 _26957_ (.A(_03943_),
    .B1(_03657_),
    .B2(_06386_),
    .ZN(_03944_));
 AND2_X4 _26958_ (.A1(_03942_),
    .A2(_03944_),
    .ZN(_03945_));
 AOI221_X2 _26959_ (.A(_03619_),
    .B1(_03709_),
    .B2(_03797_),
    .C1(_03941_),
    .C2(_03945_),
    .ZN(_03946_));
 AOI21_X2 _26960_ (.A(_15204_),
    .B1(_03663_),
    .B2(_03666_),
    .ZN(_03947_));
 AOI211_X2 _26961_ (.A(_03622_),
    .B(_03947_),
    .C1(_03797_),
    .C2(_03675_),
    .ZN(_03948_));
 OAI21_X2 _26962_ (.A(_03762_),
    .B1(_03946_),
    .B2(_03948_),
    .ZN(_03949_));
 NAND3_X1 _26963_ (.A1(_03913_),
    .A2(_03861_),
    .A3(_03824_),
    .ZN(_03950_));
 AOI21_X1 _26964_ (.A(_03707_),
    .B1(_03757_),
    .B2(_03732_),
    .ZN(_03951_));
 AOI21_X1 _26965_ (.A(_03714_),
    .B1(_03950_),
    .B2(_03951_),
    .ZN(_03952_));
 INV_X1 _26966_ (.A(_15215_),
    .ZN(_03953_));
 OAI221_X1 _26967_ (.A(_03632_),
    .B1(_03802_),
    .B2(_03764_),
    .C1(_03727_),
    .C2(_03953_),
    .ZN(_03954_));
 NOR3_X1 _26968_ (.A1(net153),
    .A2(_03727_),
    .A3(_03854_),
    .ZN(_03955_));
 OAI21_X1 _26969_ (.A(_03708_),
    .B1(_03677_),
    .B2(_15224_),
    .ZN(_03956_));
 OAI21_X1 _26970_ (.A(_03954_),
    .B1(_03955_),
    .B2(_03956_),
    .ZN(_03957_));
 AOI221_X2 _26971_ (.A(_03821_),
    .B1(_03949_),
    .B2(_03952_),
    .C1(_03957_),
    .C2(_03715_),
    .ZN(_03958_));
 OR2_X2 _26972_ (.A1(_03698_),
    .A2(_03958_),
    .ZN(_03959_));
 AOI21_X1 _26973_ (.A(_03720_),
    .B1(_03728_),
    .B2(_03846_),
    .ZN(_03960_));
 AOI21_X4 _26974_ (.A(_15210_),
    .B1(_03664_),
    .B2(_03667_),
    .ZN(_03961_));
 NOR3_X1 _26975_ (.A1(_03845_),
    .A2(_03889_),
    .A3(_03961_),
    .ZN(_03962_));
 NOR3_X1 _26976_ (.A1(_15206_),
    .A2(_03794_),
    .A3(_03795_),
    .ZN(_03963_));
 NOR3_X1 _26977_ (.A1(_03720_),
    .A2(_03847_),
    .A3(_03963_),
    .ZN(_03964_));
 NOR2_X1 _26978_ (.A1(_03716_),
    .A2(_03727_),
    .ZN(_03965_));
 NOR3_X1 _26979_ (.A1(_03687_),
    .A2(_03965_),
    .A3(_03961_),
    .ZN(_03966_));
 OAI33_X1 _26980_ (.A1(_03822_),
    .A2(_03960_),
    .A3(_03962_),
    .B1(_03964_),
    .B2(_03966_),
    .B3(_03747_),
    .ZN(_03967_));
 OR3_X1 _26981_ (.A1(_03760_),
    .A2(_03819_),
    .A3(_03967_),
    .ZN(_03968_));
 NAND2_X1 _26982_ (.A1(_03861_),
    .A2(_03897_),
    .ZN(_03969_));
 AOI221_X2 _26983_ (.A(_03715_),
    .B1(_03728_),
    .B2(_03896_),
    .C1(_03969_),
    .C2(_15212_),
    .ZN(_03970_));
 INV_X2 _26984_ (.A(_15206_),
    .ZN(_03971_));
 NOR2_X2 _26985_ (.A1(_03971_),
    .A2(_03676_),
    .ZN(_03972_));
 NOR3_X1 _26986_ (.A1(_15219_),
    .A2(_03972_),
    .A3(_03965_),
    .ZN(_03973_));
 NOR3_X1 _26987_ (.A1(_03820_),
    .A2(_03914_),
    .A3(_03973_),
    .ZN(_03974_));
 NOR3_X1 _26988_ (.A1(_03865_),
    .A2(_03970_),
    .A3(_03974_),
    .ZN(_03975_));
 OAI221_X2 _26989_ (.A(_03919_),
    .B1(_03938_),
    .B2(_03959_),
    .C1(_03968_),
    .C2(_03975_),
    .ZN(_00130_));
 OAI221_X1 _26990_ (.A(_03772_),
    .B1(_03671_),
    .B2(_03766_),
    .C1(_03802_),
    .C2(_03738_),
    .ZN(_03976_));
 NAND2_X4 _26991_ (.A1(_03605_),
    .A2(_03622_),
    .ZN(_03977_));
 OAI22_X1 _26992_ (.A1(_03894_),
    .A2(_03977_),
    .B1(_03805_),
    .B2(_15203_),
    .ZN(_03978_));
 AOI21_X1 _26993_ (.A(_03976_),
    .B1(_03978_),
    .B2(net157),
    .ZN(_03979_));
 NAND3_X1 _26994_ (.A1(_03603_),
    .A2(_03664_),
    .A3(_03667_),
    .ZN(_03980_));
 NOR2_X1 _26995_ (.A1(_03586_),
    .A2(_03980_),
    .ZN(_03981_));
 OAI21_X1 _26996_ (.A(_03762_),
    .B1(_03802_),
    .B2(_03766_),
    .ZN(_03982_));
 NOR3_X1 _26997_ (.A1(_03903_),
    .A2(_03981_),
    .A3(_03982_),
    .ZN(_03983_));
 OR4_X2 _26998_ (.A1(_03983_),
    .A2(_03761_),
    .A3(_03979_),
    .A4(_03698_),
    .ZN(_03984_));
 AND2_X4 _26999_ (.A1(_03702_),
    .A2(net1036),
    .ZN(_03985_));
 NAND3_X2 _27000_ (.A1(_15212_),
    .A2(_03865_),
    .A3(_03985_),
    .ZN(_03986_));
 NOR2_X1 _27001_ (.A1(_03661_),
    .A2(_03972_),
    .ZN(_03987_));
 AOI21_X1 _27002_ (.A(_03701_),
    .B1(_03977_),
    .B2(_03764_),
    .ZN(_03988_));
 OAI221_X2 _27003_ (.A(_03986_),
    .B1(_03987_),
    .B2(_03778_),
    .C1(_03988_),
    .C2(_03865_),
    .ZN(_03989_));
 NAND2_X1 _27004_ (.A1(_03736_),
    .A2(_03714_),
    .ZN(_03990_));
 NOR2_X1 _27005_ (.A1(net943),
    .A2(_03623_),
    .ZN(_03991_));
 NOR2_X1 _27006_ (.A1(_03718_),
    .A2(_03991_),
    .ZN(_03992_));
 OAI21_X1 _27007_ (.A(_03992_),
    .B1(_03942_),
    .B2(_03787_),
    .ZN(_03993_));
 AOI21_X1 _27008_ (.A(_03784_),
    .B1(_03720_),
    .B2(net152),
    .ZN(_03994_));
 AOI221_X2 _27009_ (.A(_03771_),
    .B1(_03877_),
    .B2(_03993_),
    .C1(_03994_),
    .C2(_03977_),
    .ZN(_03995_));
 AOI21_X1 _27010_ (.A(_15194_),
    .B1(_03913_),
    .B2(_03683_),
    .ZN(_03996_));
 AOI221_X2 _27011_ (.A(_03996_),
    .B1(_03750_),
    .B2(net156),
    .C1(_03773_),
    .C2(_03701_),
    .ZN(_03997_));
 NOR3_X1 _27012_ (.A1(_03845_),
    .A2(_03935_),
    .A3(_03961_),
    .ZN(_03998_));
 OAI21_X4 _27013_ (.A(net1036),
    .B1(_03709_),
    .B2(_03971_),
    .ZN(_03999_));
 AOI21_X1 _27014_ (.A(_03998_),
    .B1(_03999_),
    .B2(_15212_),
    .ZN(_04000_));
 OAI221_X2 _27015_ (.A(_03698_),
    .B1(_03705_),
    .B2(_03997_),
    .C1(_04000_),
    .C2(_03747_),
    .ZN(_04001_));
 OAI221_X2 _27016_ (.A(_03984_),
    .B1(_03989_),
    .B2(_03990_),
    .C1(_03995_),
    .C2(_04001_),
    .ZN(_04002_));
 AOI21_X1 _27017_ (.A(_15212_),
    .B1(_03683_),
    .B2(_03861_),
    .ZN(_04003_));
 OAI21_X1 _27018_ (.A(_03763_),
    .B1(_03748_),
    .B2(_15203_),
    .ZN(_04004_));
 AOI221_X1 _27019_ (.A(_03801_),
    .B1(_03717_),
    .B2(_03897_),
    .C1(_03977_),
    .C2(_03668_),
    .ZN(_04005_));
 OAI221_X1 _27020_ (.A(_03761_),
    .B1(_04003_),
    .B2(_04004_),
    .C1(_04005_),
    .C2(_03865_),
    .ZN(_04006_));
 NOR2_X1 _27021_ (.A1(_03686_),
    .A2(_03889_),
    .ZN(_04007_));
 NAND2_X1 _27022_ (.A1(_03649_),
    .A2(_03742_),
    .ZN(_04008_));
 AOI221_X2 _27023_ (.A(_03864_),
    .B1(_03683_),
    .B2(_04007_),
    .C1(_04008_),
    .C2(_03793_),
    .ZN(_04009_));
 OAI33_X1 _27024_ (.A1(_03826_),
    .A2(_03778_),
    .A3(_03884_),
    .B1(_03796_),
    .B2(_03947_),
    .B3(_03924_),
    .ZN(_04010_));
 OAI21_X1 _27025_ (.A(_03820_),
    .B1(_04009_),
    .B2(_04010_),
    .ZN(_04011_));
 NAND3_X1 _27026_ (.A1(_03760_),
    .A2(_04006_),
    .A3(_04011_),
    .ZN(_04012_));
 OAI21_X1 _27027_ (.A(_03714_),
    .B1(_03794_),
    .B2(_03795_),
    .ZN(_04013_));
 NOR2_X1 _27028_ (.A1(_03767_),
    .A2(_04013_),
    .ZN(_04014_));
 AOI221_X1 _27029_ (.A(_03633_),
    .B1(_03740_),
    .B2(_04014_),
    .C1(_03701_),
    .C2(_03722_),
    .ZN(_04015_));
 NAND2_X1 _27030_ (.A1(_03845_),
    .A2(_03646_),
    .ZN(_04016_));
 MUX2_X1 _27031_ (.A(_03810_),
    .B(_04016_),
    .S(_03719_),
    .Z(_04017_));
 OAI21_X1 _27032_ (.A(_04015_),
    .B1(_04017_),
    .B2(_03738_),
    .ZN(_04018_));
 NOR2_X1 _27033_ (.A1(_03839_),
    .A2(_03758_),
    .ZN(_04019_));
 AOI221_X1 _27034_ (.A(_03705_),
    .B1(_03710_),
    .B2(_03737_),
    .C1(_04019_),
    .C2(_15206_),
    .ZN(_04020_));
 AOI21_X1 _27035_ (.A(_03624_),
    .B1(_03690_),
    .B2(_03855_),
    .ZN(_04021_));
 AOI21_X1 _27036_ (.A(_03672_),
    .B1(_03688_),
    .B2(_03689_),
    .ZN(_04022_));
 NOR3_X1 _27037_ (.A1(_03794_),
    .A2(_03795_),
    .A3(net849),
    .ZN(_04023_));
 NOR3_X1 _27038_ (.A1(_03720_),
    .A2(_04022_),
    .A3(_04023_),
    .ZN(_04024_));
 NOR3_X1 _27039_ (.A1(_03804_),
    .A2(_04021_),
    .A3(_04024_),
    .ZN(_04025_));
 NOR3_X1 _27040_ (.A1(_04025_),
    .A2(_04020_),
    .A3(_03760_),
    .ZN(_04026_));
 AOI21_X2 _27041_ (.A(_03821_),
    .B1(_04026_),
    .B2(_04018_),
    .ZN(_04027_));
 AOI22_X2 _27042_ (.A1(_03821_),
    .A2(_04002_),
    .B1(_04012_),
    .B2(_04027_),
    .ZN(_00131_));
 INV_X1 _27043_ (.A(_15208_),
    .ZN(_04028_));
 MUX2_X1 _27044_ (.A(_04028_),
    .B(_03739_),
    .S(_03677_),
    .Z(_04029_));
 NAND2_X1 _27045_ (.A1(_03771_),
    .A2(_04029_),
    .ZN(_04030_));
 NOR2_X1 _27046_ (.A1(_03730_),
    .A2(_03755_),
    .ZN(_04031_));
 AOI221_X2 _27047_ (.A(_03981_),
    .B1(_04031_),
    .B2(_03913_),
    .C1(_03773_),
    .C2(_03750_),
    .ZN(_04032_));
 OAI21_X1 _27048_ (.A(_04030_),
    .B1(_04032_),
    .B2(_03771_),
    .ZN(_04033_));
 NAND3_X1 _27049_ (.A1(_03698_),
    .A2(_03853_),
    .A3(_03818_),
    .ZN(_04034_));
 NAND3_X1 _27050_ (.A1(_03698_),
    .A2(_03763_),
    .A3(_03818_),
    .ZN(_04035_));
 NAND2_X1 _27051_ (.A1(_03586_),
    .A2(_03847_),
    .ZN(_04036_));
 AOI21_X1 _27052_ (.A(_03963_),
    .B1(_03718_),
    .B2(_03645_),
    .ZN(_04037_));
 OAI221_X1 _27053_ (.A(_04036_),
    .B1(_04037_),
    .B2(_03624_),
    .C1(_03977_),
    .C2(_03878_),
    .ZN(_04038_));
 NOR2_X1 _27054_ (.A1(_03714_),
    .A2(_03727_),
    .ZN(_04039_));
 MUX2_X1 _27055_ (.A(_03737_),
    .B(_04039_),
    .S(_03624_),
    .Z(_04040_));
 AOI21_X1 _27056_ (.A(_04038_),
    .B1(_04040_),
    .B2(net154),
    .ZN(_04041_));
 OAI22_X2 _27057_ (.A1(_04033_),
    .A2(_04034_),
    .B1(_04035_),
    .B2(_04041_),
    .ZN(_04042_));
 OAI221_X1 _27058_ (.A(_03676_),
    .B1(_03740_),
    .B2(_03707_),
    .C1(_03778_),
    .C2(_03773_),
    .ZN(_04043_));
 AOI21_X1 _27059_ (.A(_03605_),
    .B1(_03620_),
    .B2(_03632_),
    .ZN(_04044_));
 OAI21_X1 _27060_ (.A(_03977_),
    .B1(_04044_),
    .B2(net153),
    .ZN(_04045_));
 OAI21_X1 _27061_ (.A(_04043_),
    .B1(_04045_),
    .B2(_03894_),
    .ZN(_04046_));
 NAND2_X1 _27062_ (.A1(_03731_),
    .A2(_03924_),
    .ZN(_04047_));
 AOI21_X1 _27063_ (.A(_03990_),
    .B1(_04047_),
    .B2(net153),
    .ZN(_04048_));
 NOR2_X1 _27064_ (.A1(_03736_),
    .A2(_03646_),
    .ZN(_04049_));
 OAI221_X2 _27065_ (.A(_03708_),
    .B1(_03868_),
    .B2(_03891_),
    .C1(_03869_),
    .C2(_03913_),
    .ZN(_04050_));
 OAI22_X1 _27066_ (.A1(net152),
    .A2(_03802_),
    .B1(_03847_),
    .B2(_03647_),
    .ZN(_04051_));
 OAI21_X2 _27067_ (.A(_04050_),
    .B1(_04051_),
    .B2(_03762_),
    .ZN(_04052_));
 AOI221_X2 _27068_ (.A(_03818_),
    .B1(_04046_),
    .B2(_04048_),
    .C1(_04049_),
    .C2(_04052_),
    .ZN(_04053_));
 NOR2_X2 _27069_ (.A1(_03971_),
    .A2(_03709_),
    .ZN(_04054_));
 AOI21_X1 _27070_ (.A(_04054_),
    .B1(_03886_),
    .B2(_03623_),
    .ZN(_04055_));
 NAND3_X1 _27071_ (.A1(_03621_),
    .A2(_03824_),
    .A3(_03871_),
    .ZN(_04056_));
 NOR2_X1 _27072_ (.A1(_03708_),
    .A2(_03710_),
    .ZN(_04057_));
 AOI221_X2 _27073_ (.A(_03697_),
    .B1(_03762_),
    .B2(_04055_),
    .C1(_04056_),
    .C2(_04057_),
    .ZN(_04058_));
 NOR2_X1 _27074_ (.A1(_03913_),
    .A2(_03632_),
    .ZN(_04059_));
 NOR2_X1 _27075_ (.A1(_03700_),
    .A2(_03620_),
    .ZN(_04060_));
 OAI21_X1 _27076_ (.A(_03718_),
    .B1(_03929_),
    .B2(_04060_),
    .ZN(_04061_));
 NOR2_X1 _27077_ (.A1(_03708_),
    .A2(_03711_),
    .ZN(_04062_));
 AOI221_X1 _27078_ (.A(_03736_),
    .B1(_04059_),
    .B2(_03887_),
    .C1(_04061_),
    .C2(_04062_),
    .ZN(_04063_));
 OAI21_X1 _27079_ (.A(_03820_),
    .B1(_04058_),
    .B2(_04063_),
    .ZN(_04064_));
 NAND2_X1 _27080_ (.A1(_03760_),
    .A2(_03819_),
    .ZN(_04065_));
 INV_X1 _27081_ (.A(_04065_),
    .ZN(_04066_));
 NOR2_X1 _27082_ (.A1(_03779_),
    .A2(_03933_),
    .ZN(_04067_));
 OAI221_X1 _27083_ (.A(_03623_),
    .B1(_03709_),
    .B2(_03773_),
    .C1(_03897_),
    .C2(net513),
    .ZN(_04068_));
 OAI21_X1 _27084_ (.A(_03702_),
    .B1(_03676_),
    .B2(_03732_),
    .ZN(_04069_));
 OAI21_X1 _27085_ (.A(_04068_),
    .B1(_04069_),
    .B2(_03913_),
    .ZN(_04070_));
 AOI221_X1 _27086_ (.A(_03908_),
    .B1(_04067_),
    .B2(_03912_),
    .C1(_04070_),
    .C2(_03772_),
    .ZN(_04071_));
 NAND2_X2 _27087_ (.A1(net156),
    .A2(_03730_),
    .ZN(_04072_));
 NOR2_X1 _27088_ (.A1(_03620_),
    .A2(_03961_),
    .ZN(_04073_));
 AOI221_X2 _27089_ (.A(_03704_),
    .B1(_04072_),
    .B2(_04073_),
    .C1(_03999_),
    .C2(_03621_),
    .ZN(_04074_));
 NAND2_X1 _27090_ (.A1(_03971_),
    .A2(_03687_),
    .ZN(_04075_));
 NAND3_X1 _27091_ (.A1(_03787_),
    .A2(_03823_),
    .A3(_03850_),
    .ZN(_04076_));
 AOI21_X1 _27092_ (.A(_03747_),
    .B1(_04075_),
    .B2(_04076_),
    .ZN(_04077_));
 OR3_X2 _27093_ (.A1(_04071_),
    .A2(_04074_),
    .A3(_04077_),
    .ZN(_04078_));
 AOI221_X2 _27094_ (.A(_04042_),
    .B1(_04064_),
    .B2(_04053_),
    .C1(_04078_),
    .C2(_04066_),
    .ZN(_00132_));
 NAND3_X1 _27095_ (.A1(net850),
    .A2(_03719_),
    .A3(_03710_),
    .ZN(_04079_));
 OAI21_X1 _27096_ (.A(_04079_),
    .B1(_03719_),
    .B2(_03766_),
    .ZN(_04080_));
 OAI22_X1 _27097_ (.A1(_03691_),
    .A2(_03872_),
    .B1(_03942_),
    .B2(_03671_),
    .ZN(_04081_));
 OAI221_X2 _27098_ (.A(_03819_),
    .B1(_03804_),
    .B2(_04080_),
    .C1(_04081_),
    .C2(_03705_),
    .ZN(_04082_));
 AOI211_X2 _27099_ (.A(_03913_),
    .B(_03961_),
    .C1(_03677_),
    .C2(net187),
    .ZN(_04083_));
 NOR3_X4 _27100_ (.A1(_03792_),
    .A2(_15219_),
    .A3(_03884_),
    .ZN(_04084_));
 NOR3_X4 _27101_ (.A1(_03820_),
    .A2(_04083_),
    .A3(_04084_),
    .ZN(_04085_));
 NAND2_X1 _27102_ (.A1(_03732_),
    .A2(_03621_),
    .ZN(_04086_));
 AOI22_X1 _27103_ (.A1(_03649_),
    .A2(_03758_),
    .B1(_04086_),
    .B2(_03719_),
    .ZN(_04087_));
 OAI21_X1 _27104_ (.A(_03865_),
    .B1(_03761_),
    .B2(_04087_),
    .ZN(_04088_));
 NOR2_X2 _27105_ (.A1(_04085_),
    .A2(_04088_),
    .ZN(_04089_));
 AOI21_X1 _27106_ (.A(_03913_),
    .B1(_03727_),
    .B2(_03971_),
    .ZN(_04090_));
 AOI221_X2 _27107_ (.A(_03747_),
    .B1(_04072_),
    .B2(_04090_),
    .C1(_03885_),
    .C2(_03683_),
    .ZN(_04091_));
 AOI22_X1 _27108_ (.A1(_15194_),
    .A2(_03691_),
    .B1(_03710_),
    .B2(_03737_),
    .ZN(_04092_));
 OAI21_X1 _27109_ (.A(_03698_),
    .B1(_03705_),
    .B2(_04092_),
    .ZN(_04093_));
 AOI21_X1 _27110_ (.A(_03894_),
    .B1(_03977_),
    .B2(_04086_),
    .ZN(_04094_));
 NOR4_X1 _27111_ (.A1(_04094_),
    .A2(_03771_),
    .A3(_03711_),
    .A4(_03763_),
    .ZN(_04095_));
 AND3_X1 _27112_ (.A1(_03624_),
    .A2(_03737_),
    .A3(_03797_),
    .ZN(_04096_));
 NOR3_X1 _27113_ (.A1(_03822_),
    .A2(_04083_),
    .A3(_04096_),
    .ZN(_04097_));
 NOR4_X2 _27114_ (.A1(_04097_),
    .A2(_04093_),
    .A3(_04095_),
    .A4(_04091_),
    .ZN(_04098_));
 OAI22_X2 _27115_ (.A1(_04089_),
    .A2(_04082_),
    .B1(_04098_),
    .B2(_03918_),
    .ZN(_04099_));
 AOI221_X1 _27116_ (.A(_03747_),
    .B1(_03894_),
    .B2(_03732_),
    .C1(_03722_),
    .C2(_03701_),
    .ZN(_04100_));
 OAI21_X1 _27117_ (.A(_04100_),
    .B1(_03991_),
    .B2(_03765_),
    .ZN(_04101_));
 NOR2_X1 _27118_ (.A1(_03698_),
    .A2(_03819_),
    .ZN(_04102_));
 AOI22_X1 _27119_ (.A1(net195),
    .A2(_03730_),
    .B1(_03850_),
    .B2(_15212_),
    .ZN(_04103_));
 OR2_X1 _27120_ (.A1(_03822_),
    .A2(_04103_),
    .ZN(_04104_));
 NAND3_X1 _27121_ (.A1(_04101_),
    .A2(_04102_),
    .A3(_04104_),
    .ZN(_04105_));
 OR3_X1 _27122_ (.A1(_15219_),
    .A2(_03889_),
    .A3(_03755_),
    .ZN(_04106_));
 AOI21_X1 _27123_ (.A(_03761_),
    .B1(_03669_),
    .B2(_04106_),
    .ZN(_04107_));
 OAI22_X1 _27124_ (.A1(_15194_),
    .A2(_03805_),
    .B1(_03999_),
    .B2(_15219_),
    .ZN(_04108_));
 OAI21_X1 _27125_ (.A(_03853_),
    .B1(_03820_),
    .B2(_04108_),
    .ZN(_04109_));
 NOR2_X1 _27126_ (.A1(_04107_),
    .A2(_04109_),
    .ZN(_04110_));
 AOI21_X1 _27127_ (.A(_03796_),
    .B1(_03719_),
    .B2(_15210_),
    .ZN(_04111_));
 OAI221_X1 _27128_ (.A(_03633_),
    .B1(_03671_),
    .B2(_03738_),
    .C1(_04111_),
    .C2(_03845_),
    .ZN(_04112_));
 OAI21_X1 _27129_ (.A(_03763_),
    .B1(_03748_),
    .B2(net850),
    .ZN(_04113_));
 NAND2_X1 _27130_ (.A1(_03722_),
    .A2(_03719_),
    .ZN(_04114_));
 AOI21_X1 _27131_ (.A(_15212_),
    .B1(_03823_),
    .B2(_04114_),
    .ZN(_04115_));
 OAI21_X1 _27132_ (.A(_04112_),
    .B1(_04113_),
    .B2(_04115_),
    .ZN(_04116_));
 NAND3_X1 _27133_ (.A1(net154),
    .A2(_03633_),
    .A3(_03802_),
    .ZN(_04117_));
 OAI21_X1 _27134_ (.A(net157),
    .B1(_03762_),
    .B2(_03894_),
    .ZN(_04118_));
 AOI21_X1 _27135_ (.A(_04118_),
    .B1(_03808_),
    .B2(_03845_),
    .ZN(_04119_));
 NOR2_X1 _27136_ (.A1(_03632_),
    .A2(_03676_),
    .ZN(_04120_));
 OAI21_X1 _27137_ (.A(_15203_),
    .B1(_04120_),
    .B2(net157),
    .ZN(_04121_));
 AOI22_X1 _27138_ (.A1(_15194_),
    .A2(_03839_),
    .B1(_03758_),
    .B2(net187),
    .ZN(_04122_));
 OAI221_X1 _27139_ (.A(_04117_),
    .B1(_04119_),
    .B2(_04121_),
    .C1(_04122_),
    .C2(_03853_),
    .ZN(_04123_));
 MUX2_X1 _27140_ (.A(_04116_),
    .B(_04123_),
    .S(_03820_),
    .Z(_04124_));
 OAI221_X2 _27141_ (.A(_04099_),
    .B1(_04105_),
    .B2(_04110_),
    .C1(_04065_),
    .C2(_04124_),
    .ZN(_00133_));
 OAI21_X1 _27142_ (.A(_03687_),
    .B1(_03891_),
    .B2(_04054_),
    .ZN(_04125_));
 AOI21_X1 _27143_ (.A(_03772_),
    .B1(_03758_),
    .B2(_03722_),
    .ZN(_04126_));
 NAND3_X1 _27144_ (.A1(_03681_),
    .A2(_03682_),
    .A3(_03623_),
    .ZN(_04127_));
 AND3_X1 _27145_ (.A1(_03676_),
    .A2(_03797_),
    .A3(_04127_),
    .ZN(_04128_));
 NOR3_X1 _27146_ (.A1(_15213_),
    .A2(_15222_),
    .A3(_03677_),
    .ZN(_04129_));
 OR2_X1 _27147_ (.A1(_04128_),
    .A2(_04129_),
    .ZN(_04130_));
 AOI221_X1 _27148_ (.A(_03818_),
    .B1(_04125_),
    .B2(_04126_),
    .C1(_04130_),
    .C2(_03853_),
    .ZN(_04131_));
 NOR2_X1 _27149_ (.A1(_03686_),
    .A2(_03755_),
    .ZN(_04132_));
 AOI221_X2 _27150_ (.A(_03704_),
    .B1(_04072_),
    .B2(_04132_),
    .C1(_03985_),
    .C2(_03687_),
    .ZN(_04133_));
 AOI221_X2 _27151_ (.A(_03894_),
    .B1(_03684_),
    .B2(net156),
    .C1(_03624_),
    .C2(net155),
    .ZN(_04134_));
 OAI21_X1 _27152_ (.A(_03763_),
    .B1(_03719_),
    .B2(_15215_),
    .ZN(_04135_));
 OAI21_X1 _27153_ (.A(_03818_),
    .B1(_04134_),
    .B2(_04135_),
    .ZN(_04136_));
 AOI21_X1 _27154_ (.A(_04133_),
    .B1(_04136_),
    .B2(_03820_),
    .ZN(_04137_));
 NAND4_X1 _27155_ (.A1(_03687_),
    .A2(_03772_),
    .A3(_03768_),
    .A4(_03883_),
    .ZN(_04138_));
 NAND2_X1 _27156_ (.A1(_03821_),
    .A2(_04138_),
    .ZN(_04139_));
 NOR3_X1 _27157_ (.A1(_03845_),
    .A2(_03864_),
    .A3(_03972_),
    .ZN(_04140_));
 NAND2_X1 _27158_ (.A1(_03742_),
    .A2(_03797_),
    .ZN(_04141_));
 AOI21_X1 _27159_ (.A(_03847_),
    .B1(_03677_),
    .B2(_15206_),
    .ZN(_04142_));
 AOI21_X1 _27160_ (.A(_04022_),
    .B1(net849),
    .B2(_03677_),
    .ZN(_04143_));
 MUX2_X1 _27161_ (.A(_04142_),
    .B(_04143_),
    .S(_03787_),
    .Z(_04144_));
 AOI221_X2 _27162_ (.A(_04139_),
    .B1(_04140_),
    .B2(_04141_),
    .C1(_03865_),
    .C2(_04144_),
    .ZN(_04145_));
 NOR2_X1 _27163_ (.A1(_03722_),
    .A2(_03732_),
    .ZN(_04146_));
 AOI21_X1 _27164_ (.A(_03621_),
    .B1(_03718_),
    .B2(_04146_),
    .ZN(_04147_));
 NOR2_X1 _27165_ (.A1(_03935_),
    .A2(_03792_),
    .ZN(_04148_));
 AOI221_X2 _27166_ (.A(_03864_),
    .B1(_04147_),
    .B2(_04072_),
    .C1(_04148_),
    .C2(_03720_),
    .ZN(_04149_));
 AOI21_X1 _27167_ (.A(_03719_),
    .B1(_03977_),
    .B2(net195),
    .ZN(_04150_));
 OAI21_X1 _27168_ (.A(_03763_),
    .B1(_03802_),
    .B2(net187),
    .ZN(_04151_));
 OAI21_X1 _27169_ (.A(_03819_),
    .B1(_04150_),
    .B2(_04151_),
    .ZN(_04152_));
 OAI21_X1 _27170_ (.A(_03761_),
    .B1(_04149_),
    .B2(_04152_),
    .ZN(_04153_));
 OAI221_X1 _27171_ (.A(_03760_),
    .B1(_04137_),
    .B2(_04131_),
    .C1(_04145_),
    .C2(_04153_),
    .ZN(_04154_));
 NOR2_X1 _27172_ (.A1(_03714_),
    .A2(_03818_),
    .ZN(_04155_));
 NAND2_X1 _27173_ (.A1(_03772_),
    .A2(_03894_),
    .ZN(_04156_));
 AOI22_X2 _27174_ (.A1(_03772_),
    .A2(_03786_),
    .B1(_03686_),
    .B2(_03961_),
    .ZN(_04157_));
 OAI221_X1 _27175_ (.A(_04155_),
    .B1(_04156_),
    .B2(_03977_),
    .C1(_04157_),
    .C2(net154),
    .ZN(_04158_));
 AOI21_X1 _27176_ (.A(_03826_),
    .B1(_03830_),
    .B2(net153),
    .ZN(_04159_));
 OAI221_X2 _27177_ (.A(_03786_),
    .B1(_04159_),
    .B2(net152),
    .C1(net157),
    .C2(_03980_),
    .ZN(_04160_));
 AOI21_X1 _27178_ (.A(_04158_),
    .B1(_04160_),
    .B2(_03763_),
    .ZN(_04161_));
 AND2_X1 _27179_ (.A1(_03686_),
    .A2(_03784_),
    .ZN(_04162_));
 OAI21_X1 _27180_ (.A(_04162_),
    .B1(_03999_),
    .B2(_03864_),
    .ZN(_04163_));
 MUX2_X1 _27181_ (.A(net512),
    .B(_03730_),
    .S(_03632_),
    .Z(_04164_));
 AOI221_X2 _27182_ (.A(_03817_),
    .B1(_04120_),
    .B2(_15203_),
    .C1(_04164_),
    .C2(_03647_),
    .ZN(_04165_));
 AOI21_X1 _27183_ (.A(_03771_),
    .B1(_04163_),
    .B2(_04165_),
    .ZN(_04166_));
 NAND2_X1 _27184_ (.A1(net154),
    .A2(_03701_),
    .ZN(_04167_));
 AOI22_X1 _27185_ (.A1(_03743_),
    .A2(_03750_),
    .B1(_03758_),
    .B2(_03971_),
    .ZN(_04168_));
 NAND3_X1 _27186_ (.A1(_03864_),
    .A2(_04167_),
    .A3(_04168_),
    .ZN(_04169_));
 OAI211_X2 _27187_ (.A(_03818_),
    .B(_04169_),
    .C1(_03916_),
    .C2(_03864_),
    .ZN(_04170_));
 NOR2_X1 _27188_ (.A1(_03761_),
    .A2(_03821_),
    .ZN(_04171_));
 NAND2_X1 _27189_ (.A1(_15214_),
    .A2(_03742_),
    .ZN(_04172_));
 OAI221_X1 _27190_ (.A(_03740_),
    .B1(_03795_),
    .B2(_03794_),
    .C1(_03971_),
    .C2(_03624_),
    .ZN(_04173_));
 AOI21_X1 _27191_ (.A(_03864_),
    .B1(_04172_),
    .B2(_04173_),
    .ZN(_04174_));
 AOI21_X1 _27192_ (.A(_04021_),
    .B1(_03701_),
    .B2(net155),
    .ZN(_04175_));
 AOI21_X1 _27193_ (.A(_04174_),
    .B1(_04175_),
    .B2(_03763_),
    .ZN(_04176_));
 AOI221_X1 _27194_ (.A(_04161_),
    .B1(_04166_),
    .B2(_04170_),
    .C1(_04171_),
    .C2(_04176_),
    .ZN(_04177_));
 OAI21_X1 _27195_ (.A(_04154_),
    .B1(_04177_),
    .B2(_03760_),
    .ZN(_00134_));
 OAI21_X1 _27196_ (.A(_03787_),
    .B1(_04013_),
    .B2(_03722_),
    .ZN(_04178_));
 NAND2_X1 _27197_ (.A1(_15203_),
    .A2(_03646_),
    .ZN(_04179_));
 OAI21_X1 _27198_ (.A(_03878_),
    .B1(_04179_),
    .B2(_03894_),
    .ZN(_04180_));
 AOI221_X2 _27199_ (.A(_04178_),
    .B1(_04180_),
    .B2(net195),
    .C1(_04039_),
    .C2(net187),
    .ZN(_04181_));
 MUX2_X1 _27200_ (.A(net745),
    .B(_03738_),
    .S(_04039_),
    .Z(_04182_));
 OAI21_X1 _27201_ (.A(_03853_),
    .B1(_04182_),
    .B2(_15219_),
    .ZN(_04183_));
 NAND3_X1 _27202_ (.A1(_03845_),
    .A2(_03941_),
    .A3(_03945_),
    .ZN(_04184_));
 OAI221_X1 _27203_ (.A(_04184_),
    .B1(_04142_),
    .B2(_03845_),
    .C1(net195),
    .C2(_03742_),
    .ZN(_04185_));
 NOR2_X1 _27204_ (.A1(_03733_),
    .A2(_04128_),
    .ZN(_04186_));
 MUX2_X1 _27205_ (.A(_04185_),
    .B(_04186_),
    .S(_03761_),
    .Z(_04187_));
 OAI221_X1 _27206_ (.A(_04102_),
    .B1(_04181_),
    .B2(_04183_),
    .C1(_04187_),
    .C2(_03853_),
    .ZN(_04188_));
 AOI221_X1 _27207_ (.A(_03646_),
    .B1(_03691_),
    .B2(_03885_),
    .C1(_03969_),
    .C2(_03787_),
    .ZN(_04189_));
 MUX2_X1 _27208_ (.A(_03700_),
    .B(_03716_),
    .S(_03620_),
    .Z(_04190_));
 AOI221_X2 _27209_ (.A(_03714_),
    .B1(_03932_),
    .B2(_03977_),
    .C1(_04190_),
    .C2(_03894_),
    .ZN(_04191_));
 OR3_X1 _27210_ (.A1(_03853_),
    .A2(_04189_),
    .A3(_04191_),
    .ZN(_04192_));
 MUX2_X1 _27211_ (.A(_03674_),
    .B(_15206_),
    .S(_03913_),
    .Z(_04193_));
 MUX2_X1 _27212_ (.A(_15222_),
    .B(_04193_),
    .S(_03737_),
    .Z(_04194_));
 AOI22_X1 _27213_ (.A1(_03722_),
    .A2(_03720_),
    .B1(_03688_),
    .B2(_03689_),
    .ZN(_04195_));
 AOI21_X1 _27214_ (.A(_04195_),
    .B1(_03742_),
    .B2(_15208_),
    .ZN(_04196_));
 OAI221_X1 _27215_ (.A(_03819_),
    .B1(_04194_),
    .B2(_03804_),
    .C1(_04196_),
    .C2(_03705_),
    .ZN(_04197_));
 INV_X1 _27216_ (.A(_04197_),
    .ZN(_04198_));
 AOI21_X2 _27217_ (.A(_03698_),
    .B1(_04198_),
    .B2(_04192_),
    .ZN(_04199_));
 AOI22_X1 _27218_ (.A1(_15219_),
    .A2(_03633_),
    .B1(_03839_),
    .B2(_03738_),
    .ZN(_04200_));
 AOI21_X1 _27219_ (.A(_03750_),
    .B1(_03742_),
    .B2(_03633_),
    .ZN(_04201_));
 OAI221_X1 _27220_ (.A(_04200_),
    .B1(_04201_),
    .B2(_03797_),
    .C1(_03912_),
    .C2(_03779_),
    .ZN(_04202_));
 AOI21_X1 _27221_ (.A(_03821_),
    .B1(_04049_),
    .B2(_04202_),
    .ZN(_04203_));
 OAI21_X1 _27222_ (.A(net154),
    .B1(_03750_),
    .B2(_03935_),
    .ZN(_04204_));
 AOI21_X1 _27223_ (.A(_03864_),
    .B1(_04036_),
    .B2(_04204_),
    .ZN(_04205_));
 AOI21_X1 _27224_ (.A(_03758_),
    .B1(_03710_),
    .B2(_03718_),
    .ZN(_04206_));
 AOI21_X1 _27225_ (.A(_03826_),
    .B1(_03701_),
    .B2(_15194_),
    .ZN(_04207_));
 OAI22_X1 _27226_ (.A1(_15195_),
    .A2(_04206_),
    .B1(_04207_),
    .B2(_03633_),
    .ZN(_04208_));
 OR4_X1 _27227_ (.A1(_03736_),
    .A2(_03761_),
    .A3(_04205_),
    .A4(_04208_),
    .ZN(_04209_));
 AOI21_X1 _27228_ (.A(_03674_),
    .B1(_03748_),
    .B2(_03805_),
    .ZN(_04210_));
 AOI221_X2 _27229_ (.A(_04210_),
    .B1(_03750_),
    .B2(_15203_),
    .C1(net152),
    .C2(_03701_),
    .ZN(_04211_));
 OAI21_X1 _27230_ (.A(_04036_),
    .B1(_03805_),
    .B2(_03797_),
    .ZN(_04212_));
 OAI221_X1 _27231_ (.A(_03771_),
    .B1(_03671_),
    .B2(_03773_),
    .C1(_03802_),
    .C2(_15203_),
    .ZN(_04213_));
 OAI221_X1 _27232_ (.A(_03865_),
    .B1(_03820_),
    .B2(_04211_),
    .C1(_04212_),
    .C2(_04213_),
    .ZN(_04214_));
 OAI21_X1 _27233_ (.A(_03787_),
    .B1(_03972_),
    .B2(_03965_),
    .ZN(_04215_));
 AOI21_X1 _27234_ (.A(_03647_),
    .B1(_03846_),
    .B2(_03883_),
    .ZN(_04216_));
 NOR2_X1 _27235_ (.A1(_03804_),
    .A2(_04216_),
    .ZN(_04217_));
 AOI22_X1 _27236_ (.A1(_03971_),
    .A2(_03758_),
    .B1(_03961_),
    .B2(_03624_),
    .ZN(_04218_));
 NAND2_X1 _27237_ (.A1(_04167_),
    .A2(_04218_),
    .ZN(_04219_));
 NOR2_X1 _27238_ (.A1(_03864_),
    .A2(_03715_),
    .ZN(_04220_));
 AOI221_X2 _27239_ (.A(_03818_),
    .B1(_04215_),
    .B2(_04217_),
    .C1(_04219_),
    .C2(_04220_),
    .ZN(_04221_));
 AOI22_X1 _27240_ (.A1(_04203_),
    .A2(_04209_),
    .B1(_04214_),
    .B2(_04221_),
    .ZN(_04222_));
 OAI21_X1 _27241_ (.A(_04188_),
    .B1(_04199_),
    .B2(_04222_),
    .ZN(_00135_));
 INV_X1 _27242_ (.A(_06341_),
    .ZN(_04223_));
 NOR2_X1 _27243_ (.A1(_04223_),
    .A2(_09179_),
    .ZN(_04224_));
 NOR2_X1 _27244_ (.A1(_06341_),
    .A2(_09179_),
    .ZN(_04225_));
 XNOR2_X2 _27245_ (.A(_12623_),
    .B(_12510_),
    .ZN(_04226_));
 XNOR2_X2 _27246_ (.A(\sa01_sr[1] ),
    .B(_09717_),
    .ZN(_04227_));
 XNOR2_X2 _27247_ (.A(_04227_),
    .B(_04226_),
    .ZN(_04228_));
 MUX2_X2 _27248_ (.A(_04224_),
    .B(_04225_),
    .S(_04228_),
    .Z(_04229_));
 OR3_X4 _27249_ (.A1(_06341_),
    .A2(_09012_),
    .A3(_00479_),
    .ZN(_04230_));
 NAND3_X2 _27250_ (.A1(_06341_),
    .A2(_09179_),
    .A3(_00479_),
    .ZN(_04231_));
 NAND2_X4 _27251_ (.A1(_04231_),
    .A2(_04230_),
    .ZN(_04232_));
 NOR2_X4 _27252_ (.A1(_04229_),
    .A2(_04232_),
    .ZN(_04233_));
 INV_X8 _27253_ (.A(net772),
    .ZN(_04234_));
 BUF_X16 _27254_ (.A(_04234_),
    .Z(_04235_));
 BUF_X32 _27255_ (.A(_04235_),
    .Z(_15232_));
 XNOR2_X1 _27256_ (.A(_09719_),
    .B(net668),
    .ZN(_04236_));
 XOR2_X2 _27257_ (.A(_09712_),
    .B(_09799_),
    .Z(_04237_));
 NAND3_X1 _27258_ (.A1(_06326_),
    .A2(_09012_),
    .A3(_04237_),
    .ZN(_04238_));
 NOR2_X1 _27259_ (.A1(_06326_),
    .A2(_09015_),
    .ZN(_04239_));
 NAND2_X1 _27260_ (.A1(net640),
    .A2(_04239_),
    .ZN(_04240_));
 AOI21_X1 _27261_ (.A(_04236_),
    .B1(_04238_),
    .B2(_04240_),
    .ZN(_04241_));
 XOR2_X1 _27262_ (.A(_09719_),
    .B(net668),
    .Z(_04242_));
 NAND2_X1 _27263_ (.A1(_04237_),
    .A2(_04239_),
    .ZN(_04243_));
 NAND3_X1 _27264_ (.A1(_06326_),
    .A2(_09194_),
    .A3(net640),
    .ZN(_04244_));
 AOI21_X1 _27265_ (.A(_04242_),
    .B1(_04243_),
    .B2(_04244_),
    .ZN(_04245_));
 INV_X1 _27266_ (.A(_06326_),
    .ZN(_04246_));
 NAND3_X1 _27267_ (.A1(_04246_),
    .A2(_09727_),
    .A3(_00480_),
    .ZN(_04247_));
 NAND2_X1 _27268_ (.A1(_06326_),
    .A2(_09028_),
    .ZN(_04248_));
 OAI21_X1 _27269_ (.A(_04247_),
    .B1(_04248_),
    .B2(_00480_),
    .ZN(_04249_));
 OR3_X4 _27270_ (.A1(_04241_),
    .A2(_04245_),
    .A3(_04249_),
    .ZN(_04250_));
 INV_X8 _27271_ (.A(_04250_),
    .ZN(_04251_));
 BUF_X4 _27272_ (.A(_04251_),
    .Z(_15235_));
 XNOR2_X1 _27273_ (.A(_09835_),
    .B(_09766_),
    .ZN(_04252_));
 NAND3_X1 _27274_ (.A1(_06356_),
    .A2(net948),
    .A3(_01593_),
    .ZN(_04253_));
 NOR2_X1 _27275_ (.A1(_06356_),
    .A2(_08970_),
    .ZN(_04254_));
 NAND2_X1 _27276_ (.A1(_12498_),
    .A2(_04254_),
    .ZN(_04255_));
 AOI21_X2 _27277_ (.A(_04252_),
    .B1(_04253_),
    .B2(_04255_),
    .ZN(_04256_));
 XNOR2_X1 _27278_ (.A(_09835_),
    .B(_09764_),
    .ZN(_04257_));
 NAND2_X1 _27279_ (.A1(_01593_),
    .A2(_04254_),
    .ZN(_04258_));
 NAND3_X1 _27280_ (.A1(_06356_),
    .A2(_09009_),
    .A3(_12498_),
    .ZN(_04259_));
 AOI21_X2 _27281_ (.A(_04257_),
    .B1(_04258_),
    .B2(_04259_),
    .ZN(_04260_));
 INV_X1 _27282_ (.A(_06356_),
    .ZN(_04261_));
 NAND3_X1 _27283_ (.A1(_04261_),
    .A2(net587),
    .A3(_00481_),
    .ZN(_04262_));
 NAND2_X1 _27284_ (.A1(_06356_),
    .A2(net587),
    .ZN(_04263_));
 OAI21_X2 _27285_ (.A(_04262_),
    .B1(_04263_),
    .B2(_00481_),
    .ZN(_04264_));
 NOR3_X4 _27286_ (.A1(_04256_),
    .A2(_04260_),
    .A3(_04264_),
    .ZN(_04265_));
 INV_X4 _27287_ (.A(_04265_),
    .ZN(_04266_));
 BUF_X4 _27288_ (.A(_04266_),
    .Z(_04267_));
 BUF_X4 _27289_ (.A(_04267_),
    .Z(_04268_));
 BUF_X4 _27290_ (.A(_04268_),
    .Z(_04269_));
 BUF_X4 _27291_ (.A(_04269_),
    .Z(_15251_));
 BUF_X16 _27292_ (.A(_04250_),
    .Z(_04270_));
 BUF_X8 _27293_ (.A(_04270_),
    .Z(_15226_));
 BUF_X4 _27294_ (.A(net1077),
    .Z(_04271_));
 BUF_X4 _27295_ (.A(_04271_),
    .Z(_04272_));
 BUF_X4 _27296_ (.A(_04272_),
    .Z(_15244_));
 XNOR2_X1 _27297_ (.A(_09798_),
    .B(_09796_),
    .ZN(_04273_));
 XNOR2_X1 _27298_ (.A(_01658_),
    .B(_04273_),
    .ZN(_04274_));
 MUX2_X2 _27299_ (.A(\text_in_r[71] ),
    .B(_04274_),
    .S(_09803_),
    .Z(_04275_));
 XNOR2_X2 _27300_ (.A(_06440_),
    .B(_04275_),
    .ZN(_04276_));
 INV_X1 _27301_ (.A(_06418_),
    .ZN(_04277_));
 XNOR2_X1 _27302_ (.A(_09872_),
    .B(_09789_),
    .ZN(_04278_));
 NOR3_X1 _27303_ (.A1(_04277_),
    .A2(_11938_),
    .A3(_04278_),
    .ZN(_04279_));
 NOR3_X1 _27304_ (.A1(_06418_),
    .A2(_11938_),
    .A3(_04278_),
    .ZN(_04280_));
 MUX2_X2 _27305_ (.A(_04279_),
    .B(_04280_),
    .S(_09816_),
    .Z(_04281_));
 XOR2_X2 _27306_ (.A(_09872_),
    .B(_09789_),
    .Z(_04282_));
 NOR3_X1 _27307_ (.A1(_06418_),
    .A2(_09102_),
    .A3(_04282_),
    .ZN(_04283_));
 NOR3_X1 _27308_ (.A1(_04277_),
    .A2(_11841_),
    .A3(_04282_),
    .ZN(_04284_));
 MUX2_X2 _27309_ (.A(_04283_),
    .B(_04284_),
    .S(_09816_),
    .Z(_04285_));
 NAND3_X1 _27310_ (.A1(_06418_),
    .A2(_09103_),
    .A3(\text_in_r[69] ),
    .ZN(_04286_));
 NAND2_X1 _27311_ (.A1(_04277_),
    .A2(_09179_),
    .ZN(_04287_));
 OAI21_X2 _27312_ (.A(_04286_),
    .B1(_04287_),
    .B2(\text_in_r[69] ),
    .ZN(_04288_));
 NOR3_X4 _27313_ (.A1(_04281_),
    .A2(_04285_),
    .A3(_04288_),
    .ZN(_04289_));
 BUF_X4 _27314_ (.A(_04289_),
    .Z(_04290_));
 NOR2_X2 _27315_ (.A1(_04276_),
    .A2(_04290_),
    .ZN(_04291_));
 XNOR2_X1 _27316_ (.A(_09788_),
    .B(_12614_),
    .ZN(_04292_));
 XNOR2_X1 _27317_ (.A(_09798_),
    .B(_04292_),
    .ZN(_04293_));
 MUX2_X2 _27318_ (.A(\text_in_r[70] ),
    .B(_04293_),
    .S(_10571_),
    .Z(_04294_));
 XNOR2_X2 _27319_ (.A(_06432_),
    .B(_04294_),
    .ZN(_04295_));
 NAND2_X1 _27320_ (.A1(_04291_),
    .A2(_04295_),
    .ZN(_04296_));
 BUF_X1 _27321_ (.A(_15228_),
    .Z(_04297_));
 INV_X2 _27322_ (.A(_04297_),
    .ZN(_04298_));
 INV_X1 _27323_ (.A(_06387_),
    .ZN(_04299_));
 NOR2_X1 _27324_ (.A1(_09194_),
    .A2(\text_in_r[67] ),
    .ZN(_04300_));
 XOR2_X2 _27325_ (.A(_09838_),
    .B(_01680_),
    .Z(_04301_));
 AOI211_X2 _27326_ (.A(_04299_),
    .B(_04300_),
    .C1(_04301_),
    .C2(_09075_),
    .ZN(_04302_));
 INV_X1 _27327_ (.A(\text_in_r[67] ),
    .ZN(_04303_));
 NOR2_X1 _27328_ (.A1(_09074_),
    .A2(_04303_),
    .ZN(_04304_));
 XNOR2_X2 _27329_ (.A(_09838_),
    .B(_01680_),
    .ZN(_04305_));
 AOI211_X2 _27330_ (.A(_06387_),
    .B(_04304_),
    .C1(_04305_),
    .C2(net1085),
    .ZN(_04306_));
 NOR3_X4 _27331_ (.A1(_04266_),
    .A2(net17),
    .A3(net11),
    .ZN(_04307_));
 NAND2_X1 _27332_ (.A1(_08995_),
    .A2(_04303_),
    .ZN(_04308_));
 OAI211_X4 _27333_ (.A(_06387_),
    .B(_04308_),
    .C1(_04305_),
    .C2(_08995_),
    .ZN(_04309_));
 BUF_X4 _27334_ (.A(_04309_),
    .Z(_04310_));
 NAND2_X1 _27335_ (.A1(_00991_),
    .A2(\text_in_r[67] ),
    .ZN(_04311_));
 OAI211_X4 _27336_ (.A(_04299_),
    .B(_04311_),
    .C1(_04301_),
    .C2(_00991_),
    .ZN(_04312_));
 BUF_X4 _27337_ (.A(_04312_),
    .Z(_04313_));
 NAND3_X4 _27338_ (.A1(_04251_),
    .A2(_04310_),
    .A3(_04313_),
    .ZN(_04314_));
 NOR2_X2 _27339_ (.A1(net17),
    .A2(net11),
    .ZN(_04315_));
 BUF_X4 _27340_ (.A(_04315_),
    .Z(_04316_));
 BUF_X4 _27341_ (.A(_04316_),
    .Z(_04317_));
 INV_X1 _27342_ (.A(net777),
    .ZN(_04318_));
 OAI21_X1 _27343_ (.A(_04314_),
    .B1(_04317_),
    .B2(_04318_),
    .ZN(_04319_));
 BUF_X4 _27344_ (.A(_04268_),
    .Z(_04320_));
 AOI22_X2 _27345_ (.A1(_04298_),
    .A2(_04307_),
    .B1(_04319_),
    .B2(_04320_),
    .ZN(_04321_));
 XNOR2_X1 _27346_ (.A(_09871_),
    .B(_01668_),
    .ZN(_04322_));
 MUX2_X2 _27347_ (.A(\text_in_r[68] ),
    .B(_04322_),
    .S(net1085),
    .Z(_04323_));
 XOR2_X2 _27348_ (.A(_06404_),
    .B(_04323_),
    .Z(_04324_));
 CLKBUF_X3 clone155 (.A(_03673_),
    .Z(net155));
 INV_X4 _27350_ (.A(net1192),
    .ZN(_04326_));
 NOR2_X4 _27351_ (.A1(_04251_),
    .A2(_04266_),
    .ZN(_04327_));
 AOI22_X4 _27352_ (.A1(_04326_),
    .A2(_04267_),
    .B1(_04327_),
    .B2(_04234_),
    .ZN(_04328_));
 NAND2_X4 _27353_ (.A1(_04309_),
    .A2(_04312_),
    .ZN(_04329_));
 BUF_X4 _27354_ (.A(_04329_),
    .Z(_04330_));
 AOI21_X2 _27355_ (.A(_04324_),
    .B1(_04328_),
    .B2(_04330_),
    .ZN(_04331_));
 BUF_X4 _27356_ (.A(_04324_),
    .Z(_04332_));
 BUF_X4 _27357_ (.A(_04332_),
    .Z(_04333_));
 CLKBUF_X3 _27358_ (.A(_04316_),
    .Z(_04334_));
 CLKBUF_X3 _27359_ (.A(_04334_),
    .Z(_04335_));
 AOI21_X4 _27360_ (.A(net1082),
    .B1(_04309_),
    .B2(_04312_),
    .ZN(_04336_));
 BUF_X4 _27361_ (.A(_15229_),
    .Z(_04337_));
 BUF_X16 _27362_ (.A(net535),
    .Z(_04338_));
 AOI22_X2 _27363_ (.A1(_15249_),
    .A2(_04335_),
    .B1(_04336_),
    .B2(net1160),
    .ZN(_04339_));
 AOI221_X2 _27364_ (.A(_04296_),
    .B1(_04321_),
    .B2(_04331_),
    .C1(_04333_),
    .C2(_04339_),
    .ZN(_04340_));
 BUF_X4 _27365_ (.A(_04290_),
    .Z(_04341_));
 BUF_X4 _27366_ (.A(_04341_),
    .Z(_04342_));
 XNOR2_X2 _27367_ (.A(_06404_),
    .B(_04323_),
    .ZN(_04343_));
 BUF_X4 _27368_ (.A(_04343_),
    .Z(_04344_));
 CLKBUF_X3 _27369_ (.A(_04344_),
    .Z(_04345_));
 INV_X2 _27370_ (.A(_15238_),
    .ZN(_04346_));
 NOR2_X1 _27371_ (.A1(_04346_),
    .A2(_04335_),
    .ZN(_04347_));
 INV_X8 _27372_ (.A(_04337_),
    .ZN(_04348_));
 BUF_X8 _27373_ (.A(net17),
    .Z(_04349_));
 BUF_X8 _27374_ (.A(net11),
    .Z(_04350_));
 NOR3_X4 _27375_ (.A1(_04348_),
    .A2(_04349_),
    .A3(_04350_),
    .ZN(_04351_));
 NOR4_X1 _27376_ (.A1(_15251_),
    .A2(_04345_),
    .A3(_04347_),
    .A4(net780),
    .ZN(_04352_));
 XOR2_X2 _27377_ (.A(_06440_),
    .B(_04275_),
    .Z(_04353_));
 XOR2_X2 _27378_ (.A(_06432_),
    .B(_04294_),
    .Z(_04354_));
 BUF_X4 _27379_ (.A(_04354_),
    .Z(_04355_));
 NAND2_X2 _27380_ (.A1(_04353_),
    .A2(_04355_),
    .ZN(_04356_));
 NOR3_X1 _27381_ (.A1(_04342_),
    .A2(_04352_),
    .A3(_04356_),
    .ZN(_04357_));
 NAND3_X2 _27382_ (.A1(_04270_),
    .A2(_04310_),
    .A3(_04313_),
    .ZN(_04358_));
 NOR2_X2 _27383_ (.A1(_04324_),
    .A2(_04358_),
    .ZN(_04359_));
 BUF_X4 _27384_ (.A(_04317_),
    .Z(_04360_));
 CLKBUF_X3 _27385_ (.A(_04360_),
    .Z(_04361_));
 CLKBUF_X3 _27386_ (.A(net1197),
    .Z(_04362_));
 OAI21_X1 _27387_ (.A(_15251_),
    .B1(_04361_),
    .B2(_04362_),
    .ZN(_04363_));
 OAI21_X2 _27388_ (.A(_04251_),
    .B1(net767),
    .B2(net493),
    .ZN(_04364_));
 AOI21_X1 _27389_ (.A(_04333_),
    .B1(_04364_),
    .B2(_04361_),
    .ZN(_04365_));
 OAI22_X2 _27390_ (.A1(_04359_),
    .A2(_04363_),
    .B1(_04365_),
    .B2(_15251_),
    .ZN(_04366_));
 AOI21_X2 _27391_ (.A(_04340_),
    .B1(_04357_),
    .B2(_04366_),
    .ZN(_04367_));
 NAND2_X1 _27392_ (.A1(_04295_),
    .A2(_04344_),
    .ZN(_04368_));
 BUF_X8 clone195 (.A(net850),
    .Z(net195));
 INV_X4 _27394_ (.A(_15236_),
    .ZN(_04370_));
 AOI221_X2 _27395_ (.A(_04368_),
    .B1(_04336_),
    .B2(_04370_),
    .C1(net1160),
    .C2(_04307_),
    .ZN(_04371_));
 NOR3_X4 _27396_ (.A1(net1077),
    .A2(net17),
    .A3(net11),
    .ZN(_04372_));
 AOI21_X2 _27397_ (.A(_04266_),
    .B1(_04309_),
    .B2(_04312_),
    .ZN(_04373_));
 NOR2_X2 _27398_ (.A1(_04372_),
    .A2(_04373_),
    .ZN(_04374_));
 CLKBUF_X3 _27399_ (.A(_04297_),
    .Z(_04375_));
 OAI21_X1 _27400_ (.A(_04371_),
    .B1(_04374_),
    .B2(_04375_),
    .ZN(_04376_));
 BUF_X4 _27401_ (.A(_04353_),
    .Z(_04377_));
 NOR2_X1 _27402_ (.A1(_04377_),
    .A2(_04342_),
    .ZN(_04378_));
 BUF_X4 _27403_ (.A(_04295_),
    .Z(_04379_));
 OAI22_X4 _27404_ (.A1(net491),
    .A2(net765),
    .B1(_04349_),
    .B2(_04350_),
    .ZN(_04380_));
 BUF_X4 clone196 (.A(_11308_),
    .Z(net196));
 NAND3_X4 _27406_ (.A1(_04312_),
    .A2(_04309_),
    .A3(_15242_),
    .ZN(_04382_));
 NAND3_X1 _27407_ (.A1(_15244_),
    .A2(_04380_),
    .A3(_04382_),
    .ZN(_04383_));
 NOR2_X2 _27408_ (.A1(_15235_),
    .A2(_04272_),
    .ZN(_04384_));
 OAI21_X1 _27409_ (.A(_04384_),
    .B1(_04361_),
    .B2(net1203),
    .ZN(_04385_));
 AOI21_X1 _27410_ (.A(_04379_),
    .B1(_04383_),
    .B2(_04385_),
    .ZN(_04386_));
 BUF_X8 _27411_ (.A(_04233_),
    .Z(_04387_));
 BUF_X16 _27412_ (.A(_04387_),
    .Z(_04388_));
 NAND2_X1 _27413_ (.A1(net1161),
    .A2(_04320_),
    .ZN(_04389_));
 AOI21_X4 _27414_ (.A(_04348_),
    .B1(_04309_),
    .B2(_04312_),
    .ZN(_04390_));
 BUF_X4 _27415_ (.A(net1080),
    .Z(_04391_));
 NOR2_X1 _27416_ (.A1(net535),
    .A2(_04391_),
    .ZN(_04392_));
 NAND2_X1 _27417_ (.A1(net1161),
    .A2(_04330_),
    .ZN(_04393_));
 AOI221_X2 _27418_ (.A(_04355_),
    .B1(_04389_),
    .B2(_04390_),
    .C1(_04392_),
    .C2(_04393_),
    .ZN(_04394_));
 OAI21_X1 _27419_ (.A(_04333_),
    .B1(_04386_),
    .B2(_04394_),
    .ZN(_04395_));
 BUF_X4 _27420_ (.A(_04373_),
    .Z(_04396_));
 OAI21_X4 _27421_ (.A(_04267_),
    .B1(_04349_),
    .B2(_04350_),
    .ZN(_04397_));
 NAND2_X2 _27422_ (.A1(_04251_),
    .A2(_04271_),
    .ZN(_04398_));
 BUF_X4 _27423_ (.A(_04329_),
    .Z(_04399_));
 CLKBUF_X3 _27424_ (.A(_04399_),
    .Z(_04400_));
 OAI21_X1 _27425_ (.A(_04397_),
    .B1(_04398_),
    .B2(_04400_),
    .ZN(_04401_));
 AOI222_X2 _27426_ (.A1(_04318_),
    .A2(_04396_),
    .B1(_04401_),
    .B2(net1203),
    .C1(_15226_),
    .C2(_04372_),
    .ZN(_04402_));
 NAND2_X1 _27427_ (.A1(_04354_),
    .A2(_04344_),
    .ZN(_04403_));
 OR2_X1 _27428_ (.A1(_04402_),
    .A2(_04403_),
    .ZN(_04404_));
 NAND4_X1 _27429_ (.A1(_04376_),
    .A2(_04378_),
    .A3(_04395_),
    .A4(_04404_),
    .ZN(_04405_));
 NAND2_X4 _27430_ (.A1(_04289_),
    .A2(_04343_),
    .ZN(_04406_));
 NOR2_X1 _27431_ (.A1(_04377_),
    .A2(_04406_),
    .ZN(_04407_));
 NAND2_X1 _27432_ (.A1(_06341_),
    .A2(_09195_),
    .ZN(_04408_));
 NAND2_X1 _27433_ (.A1(_04223_),
    .A2(_09195_),
    .ZN(_04409_));
 MUX2_X2 _27434_ (.A(_04408_),
    .B(_04409_),
    .S(net639),
    .Z(_04410_));
 AND2_X2 _27435_ (.A1(_04230_),
    .A2(_04231_),
    .ZN(_04411_));
 NAND4_X4 _27436_ (.A1(_04410_),
    .A2(_04411_),
    .A3(_04310_),
    .A4(_04313_),
    .ZN(_04412_));
 AOI221_X2 _27437_ (.A(_04379_),
    .B1(_04384_),
    .B2(_04412_),
    .C1(_04307_),
    .C2(_04326_),
    .ZN(_04413_));
 OAI21_X4 _27438_ (.A(net534),
    .B1(_04349_),
    .B2(_04350_),
    .ZN(_04414_));
 NAND3_X2 _27439_ (.A1(_04370_),
    .A2(_04309_),
    .A3(_04312_),
    .ZN(_04415_));
 AOI21_X1 _27440_ (.A(_15251_),
    .B1(_04414_),
    .B2(_04415_),
    .ZN(_04416_));
 AOI21_X4 _27441_ (.A(_04270_),
    .B1(_04309_),
    .B2(_04312_),
    .ZN(_04417_));
 AOI221_X1 _27442_ (.A(_04272_),
    .B1(_04334_),
    .B2(_04375_),
    .C1(_04417_),
    .C2(net916),
    .ZN(_04418_));
 NOR2_X1 _27443_ (.A1(_04416_),
    .A2(_04418_),
    .ZN(_04419_));
 NOR2_X1 _27444_ (.A1(_04355_),
    .A2(_04419_),
    .ZN(_04420_));
 OAI21_X1 _27445_ (.A(_04407_),
    .B1(_04413_),
    .B2(_04420_),
    .ZN(_04421_));
 BUF_X8 clone197 (.A(_11376_),
    .Z(net197));
 OAI21_X4 _27447_ (.A(_04270_),
    .B1(net765),
    .B2(net490),
    .ZN(_04423_));
 MUX2_X1 _27448_ (.A(net769),
    .B(_04423_),
    .S(_04329_),
    .Z(_04424_));
 AOI221_X2 _27449_ (.A(_04343_),
    .B1(_04336_),
    .B2(_04370_),
    .C1(_04424_),
    .C2(_04391_),
    .ZN(_04425_));
 OR3_X4 _27450_ (.A1(_04281_),
    .A2(_04285_),
    .A3(_04288_),
    .ZN(_04426_));
 NOR2_X1 _27451_ (.A1(_04276_),
    .A2(_04426_),
    .ZN(_04427_));
 NAND2_X1 _27452_ (.A1(_04295_),
    .A2(_04427_),
    .ZN(_04428_));
 BUF_X4 _27453_ (.A(_15238_),
    .Z(_04429_));
 MUX2_X1 _27454_ (.A(net778),
    .B(_04423_),
    .S(_04315_),
    .Z(_04430_));
 AOI221_X1 _27455_ (.A(_04324_),
    .B1(_04372_),
    .B2(_04429_),
    .C1(_04430_),
    .C2(_04271_),
    .ZN(_04431_));
 NOR3_X1 _27456_ (.A1(_04425_),
    .A2(_04428_),
    .A3(_04431_),
    .ZN(_04432_));
 BUF_X4 _27457_ (.A(_04324_),
    .Z(_04433_));
 NAND2_X1 _27458_ (.A1(_04290_),
    .A2(_04433_),
    .ZN(_04434_));
 NOR2_X1 _27459_ (.A1(_04377_),
    .A2(_04434_),
    .ZN(_04435_));
 OAI21_X4 _27460_ (.A(_04251_),
    .B1(_04349_),
    .B2(_04350_),
    .ZN(_04436_));
 NAND2_X1 _27461_ (.A1(_04354_),
    .A2(_04436_),
    .ZN(_04437_));
 OAI21_X4 _27462_ (.A(_04382_),
    .B1(_04315_),
    .B2(_04234_),
    .ZN(_04438_));
 AOI221_X2 _27463_ (.A(_04437_),
    .B1(_04267_),
    .B2(_04438_),
    .C1(net535),
    .C2(_04307_),
    .ZN(_04439_));
 NOR2_X4 _27464_ (.A1(_04270_),
    .A2(_04266_),
    .ZN(_04440_));
 AOI21_X1 _27465_ (.A(_04440_),
    .B1(_04270_),
    .B2(_04387_),
    .ZN(_04441_));
 XNOR2_X1 _27466_ (.A(_04334_),
    .B(_04441_),
    .ZN(_04442_));
 AOI21_X2 _27467_ (.A(_04439_),
    .B1(_04442_),
    .B2(_04379_),
    .ZN(_04443_));
 BUF_X4 _27468_ (.A(_04426_),
    .Z(_04444_));
 BUF_X4 _27469_ (.A(_04444_),
    .Z(_04445_));
 NOR2_X2 _27470_ (.A1(_04445_),
    .A2(_04356_),
    .ZN(_04446_));
 AOI21_X1 _27471_ (.A(net1202),
    .B1(_04310_),
    .B2(_04313_),
    .ZN(_04447_));
 NOR3_X4 _27472_ (.A1(net1192),
    .A2(_04349_),
    .A3(_04350_),
    .ZN(_04448_));
 OAI21_X1 _27473_ (.A(_04272_),
    .B1(_04447_),
    .B2(_04448_),
    .ZN(_04449_));
 OAI21_X1 _27474_ (.A(_04449_),
    .B1(_04397_),
    .B2(_04298_),
    .ZN(_04450_));
 BUF_X4 _27475_ (.A(_04271_),
    .Z(_04451_));
 NOR2_X1 _27476_ (.A1(_15236_),
    .A2(_04451_),
    .ZN(_04452_));
 OAI21_X1 _27477_ (.A(_04335_),
    .B1(_04440_),
    .B2(_04452_),
    .ZN(_04453_));
 BUF_X4 _27478_ (.A(_04267_),
    .Z(_04454_));
 AOI22_X2 _27479_ (.A1(_04338_),
    .A2(_04454_),
    .B1(_04310_),
    .B2(_04313_),
    .ZN(_04455_));
 OAI21_X4 _27480_ (.A(net1077),
    .B1(net765),
    .B2(net490),
    .ZN(_04456_));
 AOI21_X2 _27481_ (.A(_04332_),
    .B1(_04455_),
    .B2(_04456_),
    .ZN(_04457_));
 AOI22_X2 _27482_ (.A1(_04333_),
    .A2(_04450_),
    .B1(_04453_),
    .B2(_04457_),
    .ZN(_04458_));
 AOI221_X2 _27483_ (.A(_04432_),
    .B1(_04443_),
    .B2(_04435_),
    .C1(_04446_),
    .C2(_04458_),
    .ZN(_04459_));
 NAND4_X2 _27484_ (.A1(_04459_),
    .A2(_04405_),
    .A3(_04421_),
    .A4(_04367_),
    .ZN(_00136_));
 NOR2_X2 _27485_ (.A1(_04444_),
    .A2(_04344_),
    .ZN(_04460_));
 NOR2_X1 _27486_ (.A1(net773),
    .A2(_04436_),
    .ZN(_04461_));
 CLKBUF_X3 _27487_ (.A(_04454_),
    .Z(_04462_));
 AOI21_X1 _27488_ (.A(_04461_),
    .B1(_04382_),
    .B2(_04462_),
    .ZN(_04463_));
 BUF_X8 clone562 (.A(_04387_),
    .Z(net1161));
 NAND2_X1 _27490_ (.A1(net776),
    .A2(_04307_),
    .ZN(_04464_));
 AND3_X1 _27491_ (.A1(_04460_),
    .A2(_04463_),
    .A3(_04464_),
    .ZN(_04465_));
 OAI21_X1 _27492_ (.A(_04270_),
    .B1(_04372_),
    .B2(_04396_),
    .ZN(_04466_));
 NOR3_X1 _27493_ (.A1(_15226_),
    .A2(_04349_),
    .A3(_04350_),
    .ZN(_04467_));
 AOI22_X1 _27494_ (.A1(net1161),
    .A2(_04467_),
    .B1(_04336_),
    .B2(net1160),
    .ZN(_04468_));
 NAND3_X1 _27495_ (.A1(_04345_),
    .A2(_04466_),
    .A3(_04468_),
    .ZN(_04469_));
 CLKBUF_X3 _27496_ (.A(_04433_),
    .Z(_04470_));
 BUF_X4 _27497_ (.A(_04391_),
    .Z(_04471_));
 AOI21_X1 _27498_ (.A(_04298_),
    .B1(_04310_),
    .B2(_04313_),
    .ZN(_04472_));
 OAI21_X1 _27499_ (.A(_04471_),
    .B1(net779),
    .B2(_04472_),
    .ZN(_04473_));
 NAND3_X2 _27500_ (.A1(net1197),
    .A2(_04310_),
    .A3(_04313_),
    .ZN(_04474_));
 NAND3_X1 _27501_ (.A1(_04462_),
    .A2(_04436_),
    .A3(_04474_),
    .ZN(_04475_));
 NAND3_X1 _27502_ (.A1(_04470_),
    .A2(_04473_),
    .A3(_04475_),
    .ZN(_04476_));
 AOI21_X2 _27503_ (.A(_04341_),
    .B1(_04469_),
    .B2(_04476_),
    .ZN(_04477_));
 NAND2_X1 _27504_ (.A1(_04360_),
    .A2(_04364_),
    .ZN(_04478_));
 NOR3_X4 _27505_ (.A1(net534),
    .A2(net17),
    .A3(net11),
    .ZN(_04479_));
 AOI21_X1 _27506_ (.A(_04479_),
    .B1(_04330_),
    .B2(_04362_),
    .ZN(_04480_));
 MUX2_X1 _27507_ (.A(_04478_),
    .B(_04480_),
    .S(_04471_),
    .Z(_04481_));
 NOR2_X4 _27508_ (.A1(_04406_),
    .A2(_04481_),
    .ZN(_04482_));
 NOR4_X4 _27509_ (.A1(_04477_),
    .A2(_04465_),
    .A3(_04356_),
    .A4(_04482_),
    .ZN(_04483_));
 NAND2_X2 _27510_ (.A1(_04353_),
    .A2(_04379_),
    .ZN(_04484_));
 BUF_X8 _27511_ (.A(_04348_),
    .Z(_04485_));
 NOR2_X2 _27512_ (.A1(_04485_),
    .A2(_04391_),
    .ZN(_04486_));
 AOI21_X1 _27513_ (.A(_04486_),
    .B1(_04272_),
    .B2(net775),
    .ZN(_04487_));
 OAI21_X1 _27514_ (.A(_04331_),
    .B1(_04487_),
    .B2(_04400_),
    .ZN(_04488_));
 OAI22_X1 _27515_ (.A1(_04362_),
    .A2(_04397_),
    .B1(_04374_),
    .B2(net146),
    .ZN(_04489_));
 AOI21_X1 _27516_ (.A(_04290_),
    .B1(_04332_),
    .B2(_04489_),
    .ZN(_04490_));
 NAND3_X1 _27517_ (.A1(_04454_),
    .A2(_04334_),
    .A3(_04433_),
    .ZN(_04491_));
 OAI21_X1 _27518_ (.A(_04491_),
    .B1(_04393_),
    .B2(_04332_),
    .ZN(_04492_));
 NAND2_X2 _27519_ (.A1(_04267_),
    .A2(_04316_),
    .ZN(_04493_));
 OAI22_X1 _27520_ (.A1(_04320_),
    .A2(_04433_),
    .B1(_04493_),
    .B2(_15235_),
    .ZN(_04494_));
 AOI22_X2 _27521_ (.A1(_15226_),
    .A2(_04492_),
    .B1(_04494_),
    .B2(net1203),
    .ZN(_04495_));
 NAND2_X2 _27522_ (.A1(_04399_),
    .A2(_04324_),
    .ZN(_04496_));
 NAND2_X2 _27523_ (.A1(_04251_),
    .A2(_04267_),
    .ZN(_04497_));
 OAI21_X1 _27524_ (.A(_04290_),
    .B1(_04496_),
    .B2(_04497_),
    .ZN(_04498_));
 OAI21_X1 _27525_ (.A(_04334_),
    .B1(_04344_),
    .B2(_04485_),
    .ZN(_04499_));
 OAI21_X1 _27526_ (.A(_04499_),
    .B1(_04496_),
    .B2(_04362_),
    .ZN(_04500_));
 CLKBUF_X3 _27527_ (.A(_04451_),
    .Z(_04501_));
 AOI21_X1 _27528_ (.A(_04498_),
    .B1(_04500_),
    .B2(_04501_),
    .ZN(_04502_));
 AOI221_X2 _27529_ (.A(_04484_),
    .B1(_04488_),
    .B2(_04490_),
    .C1(_04495_),
    .C2(_04502_),
    .ZN(_04503_));
 OR3_X2 _27530_ (.A1(_04454_),
    .A2(_04417_),
    .A3(_04448_),
    .ZN(_04504_));
 NOR2_X1 _27531_ (.A1(net171),
    .A2(_04400_),
    .ZN(_04505_));
 NOR2_X1 _27532_ (.A1(_04375_),
    .A2(_04360_),
    .ZN(_04506_));
 OAI21_X1 _27533_ (.A(_04462_),
    .B1(_04505_),
    .B2(_04506_),
    .ZN(_04507_));
 AOI21_X2 _27534_ (.A(_04406_),
    .B1(_04504_),
    .B2(_04507_),
    .ZN(_04508_));
 NAND2_X2 _27535_ (.A1(_04276_),
    .A2(_04354_),
    .ZN(_04509_));
 NAND2_X2 _27536_ (.A1(_04426_),
    .A2(_04343_),
    .ZN(_04510_));
 OR2_X4 _27537_ (.A1(net764),
    .A2(_04461_),
    .ZN(_04511_));
 AOI221_X2 _27538_ (.A(_04510_),
    .B1(_04511_),
    .B2(_04451_),
    .C1(_15226_),
    .C2(_04336_),
    .ZN(_04512_));
 NAND2_X2 _27539_ (.A1(_04444_),
    .A2(_04433_),
    .ZN(_04513_));
 NAND2_X1 _27540_ (.A1(_04318_),
    .A2(_04399_),
    .ZN(_04514_));
 AOI21_X4 _27541_ (.A(_04250_),
    .B1(_04411_),
    .B2(_04410_),
    .ZN(_04515_));
 NAND2_X2 _27542_ (.A1(_04317_),
    .A2(_04515_),
    .ZN(_04516_));
 AOI21_X1 _27543_ (.A(_04471_),
    .B1(_04514_),
    .B2(_04516_),
    .ZN(_04517_));
 NAND2_X2 _27544_ (.A1(_04485_),
    .A2(_04316_),
    .ZN(_04518_));
 OAI21_X4 _27545_ (.A(_15242_),
    .B1(_04349_),
    .B2(_04350_),
    .ZN(_04519_));
 AND3_X4 _27546_ (.A1(_04451_),
    .A2(_04518_),
    .A3(net914),
    .ZN(_04520_));
 NOR3_X1 _27547_ (.A1(_04351_),
    .A2(_04451_),
    .A3(_04417_),
    .ZN(_04521_));
 AOI21_X2 _27548_ (.A(_04447_),
    .B1(_04317_),
    .B2(_04375_),
    .ZN(_04522_));
 NOR2_X1 _27549_ (.A1(_04320_),
    .A2(_04522_),
    .ZN(_04523_));
 OAI33_X1 _27550_ (.A1(_04513_),
    .A2(_04517_),
    .A3(_04520_),
    .B1(_04521_),
    .B2(_04523_),
    .B3(_04434_),
    .ZN(_04524_));
 NOR4_X4 _27551_ (.A1(_04512_),
    .A2(_04509_),
    .A3(_04524_),
    .A4(_04508_),
    .ZN(_04525_));
 NOR2_X2 _27552_ (.A1(_04377_),
    .A2(_04355_),
    .ZN(_04526_));
 NOR3_X1 _27553_ (.A1(_15252_),
    .A2(_04290_),
    .A3(_04400_),
    .ZN(_04527_));
 NAND2_X1 _27554_ (.A1(_04471_),
    .A2(_04515_),
    .ZN(_04528_));
 NOR2_X2 _27555_ (.A1(_04370_),
    .A2(net1077),
    .ZN(_04529_));
 NOR2_X1 _27556_ (.A1(_04335_),
    .A2(_04529_),
    .ZN(_04530_));
 AOI21_X1 _27557_ (.A(_04527_),
    .B1(_04528_),
    .B2(_04530_),
    .ZN(_04531_));
 OAI21_X2 _27558_ (.A(_04526_),
    .B1(_04531_),
    .B2(_04333_),
    .ZN(_04532_));
 NAND2_X2 _27559_ (.A1(_04270_),
    .A2(net1078),
    .ZN(_04533_));
 NAND4_X1 _27560_ (.A1(_15232_),
    .A2(_04335_),
    .A3(_04533_),
    .A4(_04497_),
    .ZN(_04534_));
 NOR2_X1 _27561_ (.A1(_04298_),
    .A2(_04451_),
    .ZN(_04535_));
 OAI21_X1 _27562_ (.A(_04400_),
    .B1(_04327_),
    .B2(_04535_),
    .ZN(_04536_));
 AOI21_X1 _27563_ (.A(_04444_),
    .B1(_04534_),
    .B2(_04536_),
    .ZN(_04537_));
 NAND3_X1 _27564_ (.A1(_04269_),
    .A2(_04380_),
    .A3(_04412_),
    .ZN(_04538_));
 AND2_X1 _27565_ (.A1(_04504_),
    .A2(_04538_),
    .ZN(_04539_));
 BUF_X4 _27566_ (.A(_04445_),
    .Z(_04540_));
 AOI21_X2 _27567_ (.A(_04537_),
    .B1(_04539_),
    .B2(_04540_),
    .ZN(_04541_));
 AOI21_X4 _27568_ (.A(_04532_),
    .B1(_04541_),
    .B2(_04333_),
    .ZN(_04542_));
 NOR4_X4 _27569_ (.A1(_04525_),
    .A2(_04503_),
    .A3(_04483_),
    .A4(_04542_),
    .ZN(_00137_));
 CLKBUF_X3 _27570_ (.A(_04344_),
    .Z(_04543_));
 NAND3_X1 _27571_ (.A1(_04272_),
    .A2(_04380_),
    .A3(_04415_),
    .ZN(_04544_));
 OAI21_X2 _27572_ (.A(_04320_),
    .B1(net803),
    .B2(_04472_),
    .ZN(_04545_));
 AOI21_X2 _27573_ (.A(_04543_),
    .B1(_04545_),
    .B2(_04544_),
    .ZN(_04546_));
 OAI21_X1 _27574_ (.A(_04456_),
    .B1(_04251_),
    .B2(_04234_),
    .ZN(_04547_));
 MUX2_X1 _27575_ (.A(_15252_),
    .B(_04547_),
    .S(_04334_),
    .Z(_04548_));
 AOI211_X2 _27576_ (.A(_04341_),
    .B(_04546_),
    .C1(_04548_),
    .C2(_04345_),
    .ZN(_04549_));
 NAND3_X1 _27577_ (.A1(_04485_),
    .A2(_04412_),
    .A3(_04456_),
    .ZN(_04550_));
 NAND3_X1 _27578_ (.A1(net171),
    .A2(_04471_),
    .A3(_04358_),
    .ZN(_04551_));
 NAND3_X1 _27579_ (.A1(_15232_),
    .A2(_04360_),
    .A3(_04533_),
    .ZN(_04552_));
 AND4_X1 _27580_ (.A1(_04470_),
    .A2(_04550_),
    .A3(_04551_),
    .A4(_04552_),
    .ZN(_04553_));
 AOI221_X1 _27581_ (.A(_04330_),
    .B1(_04327_),
    .B2(_04234_),
    .C1(_04454_),
    .C2(_04485_),
    .ZN(_04554_));
 BUF_X4 _27582_ (.A(_04360_),
    .Z(_04555_));
 INV_X1 _27583_ (.A(_15249_),
    .ZN(_04556_));
 OAI21_X1 _27584_ (.A(_04543_),
    .B1(_04555_),
    .B2(_04556_),
    .ZN(_04557_));
 OAI21_X1 _27585_ (.A(_04341_),
    .B1(_04554_),
    .B2(_04557_),
    .ZN(_04558_));
 OAI21_X1 _27586_ (.A(_04355_),
    .B1(_04553_),
    .B2(_04558_),
    .ZN(_04559_));
 NOR2_X1 _27587_ (.A1(_04270_),
    .A2(_04451_),
    .ZN(_04560_));
 NAND2_X1 _27588_ (.A1(net916),
    .A2(_04334_),
    .ZN(_04561_));
 OAI22_X2 _27589_ (.A1(_15256_),
    .A2(_04361_),
    .B1(_04560_),
    .B2(_04561_),
    .ZN(_04562_));
 NOR2_X1 _27590_ (.A1(_04391_),
    .A2(_04423_),
    .ZN(_04563_));
 CLKBUF_X3 _27591_ (.A(_04330_),
    .Z(_04564_));
 MUX2_X1 _27592_ (.A(_15247_),
    .B(_04563_),
    .S(_04564_),
    .Z(_04565_));
 OAI221_X2 _27593_ (.A(_04379_),
    .B1(_04513_),
    .B2(_04562_),
    .C1(_04565_),
    .C2(_04510_),
    .ZN(_04566_));
 NOR3_X4 _27594_ (.A1(net768),
    .A2(net591),
    .A3(_04266_),
    .ZN(_04567_));
 AOI22_X4 _27595_ (.A1(_04515_),
    .A2(_04396_),
    .B1(net1189),
    .B2(_04317_),
    .ZN(_04568_));
 AOI21_X2 _27596_ (.A(_04370_),
    .B1(_04310_),
    .B2(_04313_),
    .ZN(_04569_));
 AOI21_X1 _27597_ (.A(_04569_),
    .B1(_04515_),
    .B2(_04317_),
    .ZN(_04570_));
 OAI21_X4 _27598_ (.A(_04568_),
    .B1(_04570_),
    .B2(_04272_),
    .ZN(_04571_));
 NAND2_X1 _27599_ (.A1(_04375_),
    .A2(_04330_),
    .ZN(_04572_));
 NAND3_X1 _27600_ (.A1(_04501_),
    .A2(_04572_),
    .A3(_04518_),
    .ZN(_04573_));
 AOI21_X1 _27601_ (.A(_04470_),
    .B1(_04372_),
    .B2(_04362_),
    .ZN(_04574_));
 AOI221_X2 _27602_ (.A(_04445_),
    .B1(_04470_),
    .B2(_04571_),
    .C1(_04573_),
    .C2(_04574_),
    .ZN(_04575_));
 OAI221_X1 _27603_ (.A(_04377_),
    .B1(_04549_),
    .B2(_04559_),
    .C1(_04575_),
    .C2(_04566_),
    .ZN(_04576_));
 NOR2_X1 _27604_ (.A1(_04444_),
    .A2(_04433_),
    .ZN(_04577_));
 NOR2_X1 _27605_ (.A1(net776),
    .A2(_15244_),
    .ZN(_04578_));
 NAND3_X1 _27606_ (.A1(_04358_),
    .A2(_04436_),
    .A3(_04578_),
    .ZN(_04579_));
 INV_X1 _27607_ (.A(net830),
    .ZN(_04580_));
 NAND2_X1 _27608_ (.A1(_04580_),
    .A2(_04307_),
    .ZN(_04581_));
 NAND4_X1 _27609_ (.A1(_04577_),
    .A2(_04526_),
    .A3(_04579_),
    .A4(_04581_),
    .ZN(_04582_));
 OAI21_X1 _27610_ (.A(_04457_),
    .B1(_04328_),
    .B2(_04564_),
    .ZN(_04583_));
 NAND2_X1 _27611_ (.A1(_04444_),
    .A2(_04412_),
    .ZN(_04584_));
 NAND2_X1 _27612_ (.A1(_04314_),
    .A2(_04519_),
    .ZN(_04585_));
 AOI221_X2 _27613_ (.A(_04584_),
    .B1(_04585_),
    .B2(_04320_),
    .C1(_04362_),
    .C2(_04396_),
    .ZN(_04586_));
 CLKBUF_X3 _27614_ (.A(_04543_),
    .Z(_04587_));
 OAI22_X1 _27615_ (.A1(_04342_),
    .A2(_04583_),
    .B1(_04586_),
    .B2(_04587_),
    .ZN(_04588_));
 AOI21_X1 _27616_ (.A(_04454_),
    .B1(_04314_),
    .B2(_04414_),
    .ZN(_04589_));
 NOR3_X1 _27617_ (.A1(_15230_),
    .A2(_04349_),
    .A3(_04350_),
    .ZN(_04590_));
 NAND2_X1 _27618_ (.A1(_04454_),
    .A2(_04380_),
    .ZN(_04591_));
 OAI21_X1 _27619_ (.A(_04341_),
    .B1(_04590_),
    .B2(_04591_),
    .ZN(_04592_));
 OR2_X1 _27620_ (.A1(_04589_),
    .A2(_04592_),
    .ZN(_04593_));
 NAND3_X1 _27621_ (.A1(_04526_),
    .A2(_04588_),
    .A3(_04593_),
    .ZN(_04594_));
 NOR2_X1 _27622_ (.A1(_04377_),
    .A2(_04379_),
    .ZN(_04595_));
 AOI21_X2 _27623_ (.A(_04271_),
    .B1(_04399_),
    .B2(_04429_),
    .ZN(_04596_));
 NOR2_X1 _27624_ (.A1(_04351_),
    .A2(_04417_),
    .ZN(_04597_));
 AOI221_X2 _27625_ (.A(_04433_),
    .B1(_04518_),
    .B2(_04596_),
    .C1(_04597_),
    .C2(_04272_),
    .ZN(_04598_));
 NAND2_X2 _27626_ (.A1(_15242_),
    .A2(_04267_),
    .ZN(_04599_));
 AND2_X1 _27627_ (.A1(_04399_),
    .A2(_04599_),
    .ZN(_04600_));
 NAND2_X1 _27628_ (.A1(_04346_),
    .A2(_04271_),
    .ZN(_04601_));
 OAI21_X1 _27629_ (.A(_04601_),
    .B1(_04391_),
    .B2(net146),
    .ZN(_04602_));
 AOI221_X1 _27630_ (.A(_04344_),
    .B1(_04398_),
    .B2(_04600_),
    .C1(_04602_),
    .C2(_04360_),
    .ZN(_04603_));
 OR3_X1 _27631_ (.A1(_04540_),
    .A2(_04598_),
    .A3(_04603_),
    .ZN(_04604_));
 NAND2_X1 _27632_ (.A1(_04429_),
    .A2(_04271_),
    .ZN(_04605_));
 AOI21_X1 _27633_ (.A(_04317_),
    .B1(_04599_),
    .B2(_04605_),
    .ZN(_04606_));
 AOI221_X1 _27634_ (.A(_04606_),
    .B1(_04440_),
    .B2(_04334_),
    .C1(_04362_),
    .C2(_04372_),
    .ZN(_04607_));
 NOR3_X1 _27635_ (.A1(_15251_),
    .A2(_04347_),
    .A3(_04505_),
    .ZN(_04608_));
 OAI21_X1 _27636_ (.A(_04345_),
    .B1(_15244_),
    .B2(_04362_),
    .ZN(_04609_));
 OAI221_X1 _27637_ (.A(_04540_),
    .B1(_04587_),
    .B2(_04607_),
    .C1(_04608_),
    .C2(_04609_),
    .ZN(_04610_));
 NAND3_X1 _27638_ (.A1(_04595_),
    .A2(_04604_),
    .A3(_04610_),
    .ZN(_04611_));
 NAND4_X1 _27639_ (.A1(_04576_),
    .A2(_04582_),
    .A3(_04594_),
    .A4(_04611_),
    .ZN(_00138_));
 MUX2_X1 _27640_ (.A(_04485_),
    .B(_04429_),
    .S(_04268_),
    .Z(_04612_));
 AOI221_X1 _27641_ (.A(_04543_),
    .B1(_04372_),
    .B2(net775),
    .C1(_04612_),
    .C2(_04400_),
    .ZN(_04613_));
 AOI221_X1 _27642_ (.A(_04332_),
    .B1(_04436_),
    .B2(net171),
    .C1(_15235_),
    .C2(_04269_),
    .ZN(_04614_));
 NAND3_X4 _27643_ (.A1(net1079),
    .A2(_04309_),
    .A3(_04312_),
    .ZN(_04615_));
 OAI221_X1 _27644_ (.A(_04540_),
    .B1(_04613_),
    .B2(_04614_),
    .C1(_04615_),
    .C2(net776),
    .ZN(_04616_));
 NOR3_X1 _27645_ (.A1(_04360_),
    .A2(_04433_),
    .A3(_04392_),
    .ZN(_04617_));
 AND2_X1 _27646_ (.A1(_04528_),
    .A2(_04617_),
    .ZN(_04618_));
 NAND2_X1 _27647_ (.A1(_04316_),
    .A2(_04343_),
    .ZN(_04619_));
 NOR2_X1 _27648_ (.A1(_04370_),
    .A2(_04320_),
    .ZN(_04620_));
 NOR3_X1 _27649_ (.A1(_04619_),
    .A2(_04563_),
    .A3(_04620_),
    .ZN(_04621_));
 OAI33_X1 _27650_ (.A1(_04370_),
    .A2(_04451_),
    .A3(_04317_),
    .B1(_04358_),
    .B2(net766),
    .B3(net492),
    .ZN(_04622_));
 NOR3_X1 _27651_ (.A1(_04543_),
    .A2(_04589_),
    .A3(_04622_),
    .ZN(_04623_));
 OR4_X1 _27652_ (.A1(_04445_),
    .A2(_04618_),
    .A3(_04621_),
    .A4(_04623_),
    .ZN(_04624_));
 NAND3_X1 _27653_ (.A1(_04377_),
    .A2(_04616_),
    .A3(_04624_),
    .ZN(_04625_));
 OAI21_X1 _27654_ (.A(_04451_),
    .B1(_04334_),
    .B2(net916),
    .ZN(_04626_));
 AOI221_X1 _27655_ (.A(_04406_),
    .B1(_04626_),
    .B2(_15235_),
    .C1(_04336_),
    .C2(net1203),
    .ZN(_04627_));
 OAI21_X1 _27656_ (.A(_04627_),
    .B1(_04615_),
    .B2(_04375_),
    .ZN(_04628_));
 NOR3_X2 _27657_ (.A1(_04429_),
    .A2(_04349_),
    .A3(_04350_),
    .ZN(_04629_));
 OAI21_X2 _27658_ (.A(_04454_),
    .B1(_04569_),
    .B2(_04629_),
    .ZN(_04630_));
 NAND3_X1 _27659_ (.A1(_04543_),
    .A2(_04568_),
    .A3(_04630_),
    .ZN(_04631_));
 NAND3_X1 _27660_ (.A1(_04330_),
    .A2(_04398_),
    .A3(_04599_),
    .ZN(_04632_));
 AOI21_X1 _27661_ (.A(_04290_),
    .B1(_04332_),
    .B2(_04632_),
    .ZN(_04633_));
 AOI21_X4 _27662_ (.A(_15242_),
    .B1(_04309_),
    .B2(_04312_),
    .ZN(_04634_));
 NOR2_X1 _27663_ (.A1(_04272_),
    .A2(_04634_),
    .ZN(_04635_));
 NAND3_X2 _27664_ (.A1(_15238_),
    .A2(_04310_),
    .A3(_04313_),
    .ZN(_04636_));
 NAND2_X4 _27665_ (.A1(_04414_),
    .A2(_04636_),
    .ZN(_04637_));
 AOI22_X2 _27666_ (.A1(_04314_),
    .A2(_04635_),
    .B1(_04637_),
    .B2(_04471_),
    .ZN(_04638_));
 AOI221_X2 _27667_ (.A(_04377_),
    .B1(_04631_),
    .B2(_04633_),
    .C1(_04638_),
    .C2(_04460_),
    .ZN(_04639_));
 AOI21_X1 _27668_ (.A(_04379_),
    .B1(_04628_),
    .B2(_04639_),
    .ZN(_04640_));
 NAND3_X1 _27669_ (.A1(_04454_),
    .A2(_04382_),
    .A3(_04436_),
    .ZN(_04641_));
 AOI22_X1 _27670_ (.A1(_04485_),
    .A2(_04396_),
    .B1(_04567_),
    .B2(_04316_),
    .ZN(_04642_));
 AOI21_X1 _27671_ (.A(_04510_),
    .B1(_04641_),
    .B2(_04642_),
    .ZN(_04643_));
 OAI21_X1 _27672_ (.A(_04324_),
    .B1(_04615_),
    .B2(_04318_),
    .ZN(_04644_));
 NOR3_X1 _27673_ (.A1(_04289_),
    .A2(_04315_),
    .A3(_04529_),
    .ZN(_04645_));
 MUX2_X1 _27674_ (.A(_04372_),
    .B(_04373_),
    .S(_04289_),
    .Z(_04646_));
 AOI221_X2 _27675_ (.A(_04644_),
    .B1(_04645_),
    .B2(_04456_),
    .C1(_04348_),
    .C2(_04646_),
    .ZN(_04647_));
 AOI221_X2 _27676_ (.A(_04406_),
    .B1(_04396_),
    .B2(_04251_),
    .C1(_04429_),
    .C2(_04374_),
    .ZN(_04648_));
 NOR4_X2 _27677_ (.A1(_04377_),
    .A2(_04643_),
    .A3(_04647_),
    .A4(_04648_),
    .ZN(_04649_));
 NOR3_X1 _27678_ (.A1(_04271_),
    .A2(_04417_),
    .A3(_04479_),
    .ZN(_04650_));
 MUX2_X1 _27679_ (.A(_04297_),
    .B(_15236_),
    .S(_04329_),
    .Z(_04651_));
 AOI21_X1 _27680_ (.A(_04650_),
    .B1(_04651_),
    .B2(_04451_),
    .ZN(_04652_));
 AOI21_X1 _27681_ (.A(_04390_),
    .B1(_04316_),
    .B2(_04580_),
    .ZN(_04653_));
 AOI21_X1 _27682_ (.A(_04448_),
    .B1(_04329_),
    .B2(net772),
    .ZN(_04654_));
 MUX2_X1 _27683_ (.A(_04653_),
    .B(_04654_),
    .S(_04267_),
    .Z(_04655_));
 MUX2_X1 _27684_ (.A(_04652_),
    .B(_04655_),
    .S(_04344_),
    .Z(_04656_));
 NOR2_X1 _27685_ (.A1(net779),
    .A2(_04591_),
    .ZN(_04657_));
 NOR2_X1 _27686_ (.A1(_04360_),
    .A2(_04533_),
    .ZN(_04658_));
 AOI21_X1 _27687_ (.A(_04338_),
    .B1(_04412_),
    .B2(_04456_),
    .ZN(_04659_));
 AOI21_X1 _27688_ (.A(_04334_),
    .B1(_04423_),
    .B2(_04398_),
    .ZN(_04660_));
 OAI21_X1 _27689_ (.A(_04344_),
    .B1(_04493_),
    .B2(net916),
    .ZN(_04661_));
 OAI33_X1 _27690_ (.A1(_04345_),
    .A2(_04657_),
    .A3(_04658_),
    .B1(_04659_),
    .B2(_04660_),
    .B3(_04661_),
    .ZN(_04662_));
 AOI221_X2 _27691_ (.A(_04649_),
    .B1(_04656_),
    .B2(_04427_),
    .C1(_04662_),
    .C2(_04291_),
    .ZN(_04663_));
 AOI22_X1 _27692_ (.A1(_04625_),
    .A2(_04640_),
    .B1(_04379_),
    .B2(_04663_),
    .ZN(_00139_));
 AOI221_X1 _27693_ (.A(_04543_),
    .B1(_04514_),
    .B2(_04471_),
    .C1(_04335_),
    .C2(_04429_),
    .ZN(_04664_));
 AOI21_X1 _27694_ (.A(_04271_),
    .B1(_04316_),
    .B2(_04234_),
    .ZN(_04665_));
 AOI21_X1 _27695_ (.A(_04440_),
    .B1(_04572_),
    .B2(_04665_),
    .ZN(_04666_));
 AOI21_X1 _27696_ (.A(_04664_),
    .B1(_04666_),
    .B2(_04587_),
    .ZN(_04667_));
 NOR3_X1 _27697_ (.A1(net171),
    .A2(_04269_),
    .A3(_04332_),
    .ZN(_04668_));
 NOR2_X1 _27698_ (.A1(_04501_),
    .A2(_04543_),
    .ZN(_04669_));
 AOI21_X1 _27699_ (.A(_04668_),
    .B1(_04669_),
    .B2(_04375_),
    .ZN(_04670_));
 OAI21_X1 _27700_ (.A(_15226_),
    .B1(_04501_),
    .B2(_04470_),
    .ZN(_04671_));
 AOI21_X1 _27701_ (.A(_04440_),
    .B1(_04671_),
    .B2(net1203),
    .ZN(_04672_));
 MUX2_X1 _27702_ (.A(_04670_),
    .B(_04672_),
    .S(_04564_),
    .Z(_04673_));
 NOR2_X1 _27703_ (.A1(_04462_),
    .A2(_04543_),
    .ZN(_04674_));
 OAI21_X1 _27704_ (.A(net776),
    .B1(_04359_),
    .B2(_04674_),
    .ZN(_04675_));
 AND3_X1 _27705_ (.A1(_04291_),
    .A2(_04355_),
    .A3(_04675_),
    .ZN(_04676_));
 AOI22_X1 _27706_ (.A1(_04446_),
    .A2(_04667_),
    .B1(_04673_),
    .B2(_04676_),
    .ZN(_04677_));
 OAI21_X1 _27707_ (.A(_04474_),
    .B1(_04555_),
    .B2(_04375_),
    .ZN(_04678_));
 NAND2_X1 _27708_ (.A1(_15244_),
    .A2(_04678_),
    .ZN(_04679_));
 AOI21_X1 _27709_ (.A(_04587_),
    .B1(_04538_),
    .B2(_04679_),
    .ZN(_04680_));
 OAI21_X2 _27710_ (.A(_04345_),
    .B1(_04635_),
    .B2(_04658_),
    .ZN(_04681_));
 NAND2_X1 _27711_ (.A1(_04540_),
    .A2(_04681_),
    .ZN(_04682_));
 AOI21_X2 _27712_ (.A(_04268_),
    .B1(_04399_),
    .B2(_04326_),
    .ZN(_04683_));
 OAI21_X1 _27713_ (.A(_04314_),
    .B1(_04360_),
    .B2(_04338_),
    .ZN(_04684_));
 AOI221_X2 _27714_ (.A(_04332_),
    .B1(_04516_),
    .B2(_04683_),
    .C1(_04684_),
    .C2(_04269_),
    .ZN(_04685_));
 NAND2_X1 _27715_ (.A1(_04514_),
    .A2(_04516_),
    .ZN(_04686_));
 AOI21_X1 _27716_ (.A(_04685_),
    .B1(_04686_),
    .B2(_04669_),
    .ZN(_04687_));
 OAI221_X2 _27717_ (.A(_04595_),
    .B1(_04680_),
    .B2(_04682_),
    .C1(_04687_),
    .C2(_04540_),
    .ZN(_04688_));
 NAND2_X1 _27718_ (.A1(_04391_),
    .A2(_04399_),
    .ZN(_04689_));
 NOR2_X1 _27719_ (.A1(net770),
    .A2(_04689_),
    .ZN(_04690_));
 NOR2_X1 _27720_ (.A1(_04564_),
    .A2(_04423_),
    .ZN(_04691_));
 AOI21_X1 _27721_ (.A(_04501_),
    .B1(_04314_),
    .B2(_04572_),
    .ZN(_04692_));
 NOR4_X2 _27722_ (.A1(_04342_),
    .A2(_04690_),
    .A3(_04691_),
    .A4(_04692_),
    .ZN(_04693_));
 MUX2_X1 _27723_ (.A(_15240_),
    .B(_04486_),
    .S(_04335_),
    .Z(_04694_));
 OAI21_X1 _27724_ (.A(_04587_),
    .B1(_04694_),
    .B2(_04540_),
    .ZN(_04695_));
 NAND3_X1 _27725_ (.A1(_04444_),
    .A2(_04555_),
    .A3(_04440_),
    .ZN(_04696_));
 AOI21_X1 _27726_ (.A(_04629_),
    .B1(_04564_),
    .B2(_04341_),
    .ZN(_04697_));
 OAI221_X1 _27727_ (.A(_04696_),
    .B1(_04697_),
    .B2(_15244_),
    .C1(_04361_),
    .C2(_04423_),
    .ZN(_04698_));
 OAI21_X1 _27728_ (.A(_04397_),
    .B1(_04615_),
    .B2(_04445_),
    .ZN(_04699_));
 AOI21_X1 _27729_ (.A(_04698_),
    .B1(_04699_),
    .B2(net776),
    .ZN(_04700_));
 OAI221_X2 _27730_ (.A(_04526_),
    .B1(_04693_),
    .B2(_04695_),
    .C1(_04700_),
    .C2(_04587_),
    .ZN(_04701_));
 INV_X1 _27731_ (.A(_04484_),
    .ZN(_04702_));
 NOR2_X1 _27732_ (.A1(_04462_),
    .A2(_04634_),
    .ZN(_04703_));
 OR2_X2 _27733_ (.A1(_04329_),
    .A2(_04423_),
    .ZN(_04704_));
 AOI22_X2 _27734_ (.A1(_15251_),
    .A2(_04637_),
    .B1(_04703_),
    .B2(_04704_),
    .ZN(_04705_));
 NOR2_X1 _27735_ (.A1(_04333_),
    .A2(_04705_),
    .ZN(_04706_));
 OAI21_X1 _27736_ (.A(_04462_),
    .B1(_04555_),
    .B2(_04326_),
    .ZN(_04707_));
 OAI21_X1 _27737_ (.A(_04601_),
    .B1(_04707_),
    .B2(net780),
    .ZN(_04708_));
 OAI21_X1 _27738_ (.A(_04342_),
    .B1(_04587_),
    .B2(_04708_),
    .ZN(_04709_));
 OAI21_X2 _27739_ (.A(_04519_),
    .B1(_04330_),
    .B2(net1161),
    .ZN(_04710_));
 AOI221_X2 _27740_ (.A(_04543_),
    .B1(_04704_),
    .B2(_04683_),
    .C1(_04710_),
    .C2(_04269_),
    .ZN(_04711_));
 NOR2_X1 _27741_ (.A1(_04375_),
    .A2(_15251_),
    .ZN(_04712_));
 OAI21_X1 _27742_ (.A(_04361_),
    .B1(_04578_),
    .B2(_04712_),
    .ZN(_04713_));
 AOI21_X1 _27743_ (.A(_04711_),
    .B1(_04713_),
    .B2(_04331_),
    .ZN(_04714_));
 OAI221_X2 _27744_ (.A(_04702_),
    .B1(_04706_),
    .B2(_04709_),
    .C1(_04714_),
    .C2(_04342_),
    .ZN(_04715_));
 NAND4_X4 _27745_ (.A1(_04688_),
    .A2(_04677_),
    .A3(_04701_),
    .A4(_04715_),
    .ZN(_00140_));
 OAI21_X1 _27746_ (.A(_04519_),
    .B1(_04399_),
    .B2(_04297_),
    .ZN(_04716_));
 AOI221_X2 _27747_ (.A(_04324_),
    .B1(_04485_),
    .B2(_04307_),
    .C1(_04716_),
    .C2(_04268_),
    .ZN(_04717_));
 MUX2_X1 _27748_ (.A(net535),
    .B(net769),
    .S(_04329_),
    .Z(_04718_));
 AOI221_X1 _27749_ (.A(_04343_),
    .B1(_04396_),
    .B2(net146),
    .C1(_04718_),
    .C2(_04268_),
    .ZN(_04719_));
 NOR3_X1 _27750_ (.A1(_04717_),
    .A2(_04296_),
    .A3(_04719_),
    .ZN(_04720_));
 AOI21_X2 _27751_ (.A(net1081),
    .B1(_04329_),
    .B2(_04346_),
    .ZN(_04721_));
 AOI21_X1 _27752_ (.A(_04479_),
    .B1(_04399_),
    .B2(_04387_),
    .ZN(_04722_));
 AOI221_X2 _27753_ (.A(_04426_),
    .B1(_04704_),
    .B2(_04721_),
    .C1(_04722_),
    .C2(_04391_),
    .ZN(_04723_));
 NAND2_X1 _27754_ (.A1(_04415_),
    .A2(_04519_),
    .ZN(_04724_));
 AOI221_X2 _27755_ (.A(_04289_),
    .B1(_04364_),
    .B2(_04396_),
    .C1(_04724_),
    .C2(_04268_),
    .ZN(_04725_));
 OAI21_X1 _27756_ (.A(_04470_),
    .B1(_04725_),
    .B2(_04723_),
    .ZN(_04726_));
 AOI221_X2 _27757_ (.A(_04289_),
    .B1(_04515_),
    .B2(_04307_),
    .C1(_04326_),
    .C2(_04336_),
    .ZN(_04727_));
 OAI22_X1 _27758_ (.A1(_04316_),
    .A2(_04423_),
    .B1(_04396_),
    .B2(_04270_),
    .ZN(_04728_));
 AOI221_X2 _27759_ (.A(_04324_),
    .B1(_04466_),
    .B2(_04727_),
    .C1(_04728_),
    .C2(_04289_),
    .ZN(_04729_));
 NOR2_X2 _27760_ (.A1(_04729_),
    .A2(_04509_),
    .ZN(_04730_));
 OAI21_X1 _27761_ (.A(net776),
    .B1(_04555_),
    .B2(_04577_),
    .ZN(_04731_));
 OAI21_X1 _27762_ (.A(_04555_),
    .B1(_04577_),
    .B2(_04462_),
    .ZN(_04732_));
 NOR2_X1 _27763_ (.A1(net146),
    .A2(_04316_),
    .ZN(_04733_));
 AOI21_X1 _27764_ (.A(_15226_),
    .B1(_04733_),
    .B2(_04460_),
    .ZN(_04734_));
 NAND3_X1 _27765_ (.A1(_04731_),
    .A2(_04732_),
    .A3(_04734_),
    .ZN(_04735_));
 OAI22_X2 _27766_ (.A1(_04317_),
    .A2(_04533_),
    .B1(_04493_),
    .B2(_04370_),
    .ZN(_04736_));
 OAI21_X1 _27767_ (.A(_04317_),
    .B1(_04343_),
    .B2(_04529_),
    .ZN(_04737_));
 NAND2_X1 _27768_ (.A1(_04689_),
    .A2(_04737_),
    .ZN(_04738_));
 AOI221_X2 _27769_ (.A(_04428_),
    .B1(_04736_),
    .B2(_04433_),
    .C1(_04738_),
    .C2(net171),
    .ZN(_04739_));
 AOI221_X2 _27770_ (.A(_04720_),
    .B1(_04730_),
    .B2(_04726_),
    .C1(_04735_),
    .C2(_04739_),
    .ZN(_04740_));
 NOR2_X1 _27771_ (.A1(_04326_),
    .A2(_15244_),
    .ZN(_04741_));
 OAI221_X1 _27772_ (.A(_04333_),
    .B1(_04493_),
    .B2(net775),
    .C1(_04741_),
    .C2(_04361_),
    .ZN(_04742_));
 NAND2_X1 _27773_ (.A1(_04361_),
    .A2(net1190),
    .ZN(_04743_));
 OR3_X1 _27774_ (.A1(_04327_),
    .A2(_04380_),
    .A3(_04560_),
    .ZN(_04744_));
 NAND3_X1 _27775_ (.A1(_04345_),
    .A2(_04743_),
    .A3(_04744_),
    .ZN(_04745_));
 AOI21_X1 _27776_ (.A(_04540_),
    .B1(_04742_),
    .B2(_04745_),
    .ZN(_04746_));
 NOR3_X1 _27777_ (.A1(_04462_),
    .A2(_04390_),
    .A3(net764),
    .ZN(_04747_));
 AOI21_X1 _27778_ (.A(_04747_),
    .B1(_04724_),
    .B2(_15251_),
    .ZN(_04748_));
 NOR2_X1 _27779_ (.A1(_04513_),
    .A2(_04748_),
    .ZN(_04749_));
 AOI221_X1 _27780_ (.A(_04510_),
    .B1(_04461_),
    .B2(_04471_),
    .C1(_15236_),
    .C2(_04555_),
    .ZN(_04750_));
 NOR3_X1 _27781_ (.A1(_04746_),
    .A2(_04749_),
    .A3(_04750_),
    .ZN(_04751_));
 NAND2_X1 _27782_ (.A1(_04276_),
    .A2(_04379_),
    .ZN(_04752_));
 AOI21_X1 _27783_ (.A(_04269_),
    .B1(_04400_),
    .B2(_04362_),
    .ZN(_04753_));
 OAI21_X1 _27784_ (.A(_04445_),
    .B1(_04691_),
    .B2(_04753_),
    .ZN(_04754_));
 OAI22_X1 _27785_ (.A1(_04429_),
    .A2(_04471_),
    .B1(_04533_),
    .B2(net1161),
    .ZN(_04755_));
 NAND2_X1 _27786_ (.A1(net1202),
    .A2(_04471_),
    .ZN(_04756_));
 AOI22_X1 _27787_ (.A1(_04564_),
    .A2(_04755_),
    .B1(_04756_),
    .B2(_04448_),
    .ZN(_04757_));
 OAI21_X1 _27788_ (.A(_04754_),
    .B1(_04757_),
    .B2(_04445_),
    .ZN(_04758_));
 OAI21_X1 _27789_ (.A(_04449_),
    .B1(_04438_),
    .B2(_04501_),
    .ZN(_04759_));
 OAI22_X1 _27790_ (.A1(_15226_),
    .A2(_04493_),
    .B1(_04637_),
    .B2(_04269_),
    .ZN(_04760_));
 MUX2_X1 _27791_ (.A(_04759_),
    .B(_04760_),
    .S(_04444_),
    .Z(_04761_));
 MUX2_X1 _27792_ (.A(_04758_),
    .B(_04761_),
    .S(_04587_),
    .Z(_04762_));
 OAI221_X2 _27793_ (.A(_04740_),
    .B1(_04751_),
    .B2(_04752_),
    .C1(_04356_),
    .C2(_04762_),
    .ZN(_00141_));
 AOI22_X1 _27794_ (.A1(_04429_),
    .A2(_04320_),
    .B1(_04310_),
    .B2(_04313_),
    .ZN(_04763_));
 AOI22_X1 _27795_ (.A1(_15246_),
    .A2(_04555_),
    .B1(_04456_),
    .B2(_04763_),
    .ZN(_04764_));
 NOR2_X1 _27796_ (.A1(_04540_),
    .A2(_04764_),
    .ZN(_04765_));
 NOR3_X1 _27797_ (.A1(_04341_),
    .A2(_04564_),
    .A3(_04328_),
    .ZN(_04766_));
 OAI21_X1 _27798_ (.A(_04587_),
    .B1(_04765_),
    .B2(_04766_),
    .ZN(_04767_));
 NAND2_X1 _27799_ (.A1(_04382_),
    .A2(_04436_),
    .ZN(_04768_));
 AOI221_X1 _27800_ (.A(_04434_),
    .B1(_04768_),
    .B2(_04320_),
    .C1(_04307_),
    .C2(_04485_),
    .ZN(_04769_));
 AOI21_X1 _27801_ (.A(_04513_),
    .B1(_04630_),
    .B2(_04464_),
    .ZN(_04770_));
 NOR2_X1 _27802_ (.A1(_04769_),
    .A2(_04770_),
    .ZN(_04771_));
 AOI21_X1 _27803_ (.A(_04752_),
    .B1(_04767_),
    .B2(_04771_),
    .ZN(_04772_));
 MUX2_X1 _27804_ (.A(_04375_),
    .B(_15235_),
    .S(_04444_),
    .Z(_04773_));
 OAI21_X1 _27805_ (.A(_04636_),
    .B1(_04773_),
    .B2(_04555_),
    .ZN(_04774_));
 NAND2_X1 _27806_ (.A1(_15244_),
    .A2(_04774_),
    .ZN(_04775_));
 OAI21_X1 _27807_ (.A(_04474_),
    .B1(_04335_),
    .B2(net1160),
    .ZN(_04776_));
 AOI22_X2 _27808_ (.A1(net771),
    .A2(_04361_),
    .B1(_04776_),
    .B2(_04445_),
    .ZN(_04777_));
 OAI211_X2 _27809_ (.A(_04333_),
    .B(_04775_),
    .C1(_04777_),
    .C2(_15244_),
    .ZN(_04778_));
 AOI21_X1 _27810_ (.A(_04478_),
    .B1(_04501_),
    .B2(net776),
    .ZN(_04779_));
 OR2_X1 _27811_ (.A1(_15245_),
    .A2(_15254_),
    .ZN(_04780_));
 OAI21_X1 _27812_ (.A(_04341_),
    .B1(_04555_),
    .B2(_04780_),
    .ZN(_04781_));
 NOR3_X1 _27813_ (.A1(_04269_),
    .A2(_04590_),
    .A3(_04634_),
    .ZN(_04782_));
 AOI21_X1 _27814_ (.A(_04782_),
    .B1(_04721_),
    .B2(_04516_),
    .ZN(_04783_));
 OAI221_X1 _27815_ (.A(_04587_),
    .B1(_04779_),
    .B2(_04781_),
    .C1(_04783_),
    .C2(_04342_),
    .ZN(_04784_));
 AOI21_X1 _27816_ (.A(_04356_),
    .B1(_04778_),
    .B2(_04784_),
    .ZN(_04785_));
 OAI21_X4 _27817_ (.A(_04330_),
    .B1(_04338_),
    .B2(_04268_),
    .ZN(_04786_));
 OAI221_X2 _27818_ (.A(_04290_),
    .B1(_04786_),
    .B2(_04563_),
    .C1(_04400_),
    .C2(_15247_),
    .ZN(_04787_));
 NOR2_X1 _27819_ (.A1(_04387_),
    .A2(_04440_),
    .ZN(_04788_));
 OAI221_X1 _27820_ (.A(_04444_),
    .B1(_04400_),
    .B2(_04788_),
    .C1(_04397_),
    .C2(_15236_),
    .ZN(_04789_));
 AND3_X4 _27821_ (.A1(_04787_),
    .A2(_04470_),
    .A3(_04789_),
    .ZN(_04790_));
 NAND3_X1 _27822_ (.A1(_04501_),
    .A2(_04414_),
    .A3(_04412_),
    .ZN(_04791_));
 NAND2_X1 _27823_ (.A1(_04462_),
    .A2(_04430_),
    .ZN(_04792_));
 AOI21_X1 _27824_ (.A(_04406_),
    .B1(_04791_),
    .B2(_04792_),
    .ZN(_04793_));
 NAND2_X1 _27825_ (.A1(_04391_),
    .A2(_04704_),
    .ZN(_04794_));
 NAND3_X1 _27826_ (.A1(_04268_),
    .A2(_04314_),
    .A3(_04414_),
    .ZN(_04795_));
 AOI221_X2 _27827_ (.A(_04510_),
    .B1(_04795_),
    .B2(_04794_),
    .C1(net1191),
    .C2(_04400_),
    .ZN(_04796_));
 NOR4_X4 _27828_ (.A1(_04790_),
    .A2(_04484_),
    .A3(_04793_),
    .A4(_04796_),
    .ZN(_04797_));
 AOI22_X2 _27829_ (.A1(_04343_),
    .A2(_04497_),
    .B1(_04634_),
    .B2(_04271_),
    .ZN(_04798_));
 OAI221_X1 _27830_ (.A(_04290_),
    .B1(_04619_),
    .B2(_04398_),
    .C1(_04798_),
    .C2(_04387_),
    .ZN(_04799_));
 AOI21_X1 _27831_ (.A(_04417_),
    .B1(_04327_),
    .B2(net146),
    .ZN(_04800_));
 OAI221_X1 _27832_ (.A(_04497_),
    .B1(_04800_),
    .B2(net775),
    .C1(net916),
    .C2(_04358_),
    .ZN(_04801_));
 AOI21_X2 _27833_ (.A(_04799_),
    .B1(_04801_),
    .B2(_04470_),
    .ZN(_04802_));
 NOR2_X1 _27834_ (.A1(_04235_),
    .A2(_04344_),
    .ZN(_04803_));
 OAI21_X1 _27835_ (.A(_04320_),
    .B1(_04359_),
    .B2(_04803_),
    .ZN(_04804_));
 OAI21_X1 _27836_ (.A(_04496_),
    .B1(_04637_),
    .B2(_04433_),
    .ZN(_04805_));
 OAI221_X2 _27837_ (.A(_04804_),
    .B1(_04805_),
    .B2(_04269_),
    .C1(_15226_),
    .C2(_04496_),
    .ZN(_04806_));
 AOI211_X2 _27838_ (.A(_04509_),
    .B(_04802_),
    .C1(_04806_),
    .C2(_04445_),
    .ZN(_04807_));
 NOR4_X2 _27839_ (.A1(_04807_),
    .A2(_04785_),
    .A3(_04772_),
    .A4(_04797_),
    .ZN(_00142_));
 AOI21_X1 _27840_ (.A(_04364_),
    .B1(_04397_),
    .B2(_04619_),
    .ZN(_04808_));
 NAND4_X1 _27841_ (.A1(_04235_),
    .A2(_04360_),
    .A3(_04332_),
    .A4(_04327_),
    .ZN(_04809_));
 OAI221_X1 _27842_ (.A(_04809_),
    .B1(_04470_),
    .B2(_04501_),
    .C1(_04485_),
    .C2(_04689_),
    .ZN(_04810_));
 NOR3_X1 _27843_ (.A1(_04355_),
    .A2(_04808_),
    .A3(_04810_),
    .ZN(_04811_));
 AND2_X1 _27844_ (.A1(_04314_),
    .A2(net915),
    .ZN(_04812_));
 AOI221_X2 _27845_ (.A(_04403_),
    .B1(_04561_),
    .B2(_04596_),
    .C1(_04812_),
    .C2(_04501_),
    .ZN(_04813_));
 OAI21_X1 _27846_ (.A(_04581_),
    .B1(_04397_),
    .B2(_15235_),
    .ZN(_04814_));
 NAND2_X1 _27847_ (.A1(_04355_),
    .A2(_04470_),
    .ZN(_04815_));
 NOR2_X1 _27848_ (.A1(net1160),
    .A2(_04374_),
    .ZN(_04816_));
 NOR3_X1 _27849_ (.A1(_04814_),
    .A2(_04815_),
    .A3(_04816_),
    .ZN(_04817_));
 NOR4_X2 _27850_ (.A1(_04342_),
    .A2(_04811_),
    .A3(_04813_),
    .A4(_04817_),
    .ZN(_04818_));
 NOR2_X1 _27851_ (.A1(_04335_),
    .A2(_04423_),
    .ZN(_04819_));
 AOI21_X1 _27852_ (.A(net1203),
    .B1(_04314_),
    .B2(_04397_),
    .ZN(_04820_));
 OAI21_X1 _27853_ (.A(_04345_),
    .B1(_04819_),
    .B2(_04820_),
    .ZN(_04821_));
 AOI21_X1 _27854_ (.A(_04417_),
    .B1(_04307_),
    .B2(_15226_),
    .ZN(_04822_));
 AOI21_X1 _27855_ (.A(_04372_),
    .B1(_04396_),
    .B2(_15235_),
    .ZN(_04823_));
 OAI221_X1 _27856_ (.A(_04821_),
    .B1(_04822_),
    .B2(_04345_),
    .C1(net776),
    .C2(_04823_),
    .ZN(_04824_));
 NOR3_X1 _27857_ (.A1(_04540_),
    .A2(_04355_),
    .A3(_04824_),
    .ZN(_04825_));
 OAI221_X1 _27858_ (.A(_04333_),
    .B1(_04615_),
    .B2(_04298_),
    .C1(_04397_),
    .C2(_15235_),
    .ZN(_04826_));
 MUX2_X1 _27859_ (.A(_04564_),
    .B(_04372_),
    .S(_15235_),
    .Z(_04827_));
 AOI21_X1 _27860_ (.A(_04826_),
    .B1(_04827_),
    .B2(net1203),
    .ZN(_04828_));
 OAI221_X1 _27861_ (.A(_04345_),
    .B1(_04493_),
    .B2(_04429_),
    .C1(_04710_),
    .C2(_15251_),
    .ZN(_04829_));
 NAND3_X1 _27862_ (.A1(_04342_),
    .A2(_04355_),
    .A3(_04829_),
    .ZN(_04830_));
 OAI21_X1 _27863_ (.A(_04276_),
    .B1(_04828_),
    .B2(_04830_),
    .ZN(_04831_));
 AOI21_X1 _27864_ (.A(net1190),
    .B1(_04462_),
    .B2(_04346_),
    .ZN(_04832_));
 OAI221_X1 _27865_ (.A(_04341_),
    .B1(_04380_),
    .B2(_04384_),
    .C1(_04832_),
    .C2(_04564_),
    .ZN(_04833_));
 OAI21_X1 _27866_ (.A(_04445_),
    .B1(_04361_),
    .B2(_04362_),
    .ZN(_04834_));
 OAI21_X1 _27867_ (.A(_04833_),
    .B1(_04834_),
    .B2(_04779_),
    .ZN(_04835_));
 OAI21_X1 _27868_ (.A(_04377_),
    .B1(_04815_),
    .B2(_04835_),
    .ZN(_04836_));
 AOI221_X1 _27869_ (.A(_04289_),
    .B1(_04514_),
    .B2(_04665_),
    .C1(_04272_),
    .C2(_04298_),
    .ZN(_04837_));
 AOI22_X1 _27870_ (.A1(_15236_),
    .A2(_04335_),
    .B1(_04417_),
    .B2(_04235_),
    .ZN(_04838_));
 OAI21_X1 _27871_ (.A(_04473_),
    .B1(_04838_),
    .B2(_15244_),
    .ZN(_04839_));
 AOI21_X1 _27872_ (.A(_04837_),
    .B1(_04839_),
    .B2(_04342_),
    .ZN(_04840_));
 NOR2_X1 _27873_ (.A1(_04403_),
    .A2(_04840_),
    .ZN(_04841_));
 NAND2_X1 _27874_ (.A1(net1202),
    .A2(_04267_),
    .ZN(_04842_));
 MUX2_X1 _27875_ (.A(_15240_),
    .B(_04842_),
    .S(_04399_),
    .Z(_04843_));
 AOI21_X1 _27876_ (.A(_04332_),
    .B1(_04843_),
    .B2(_04290_),
    .ZN(_04844_));
 OAI21_X1 _27877_ (.A(_04605_),
    .B1(_04391_),
    .B2(_04338_),
    .ZN(_04845_));
 MUX2_X1 _27878_ (.A(_15254_),
    .B(_04845_),
    .S(_04330_),
    .Z(_04846_));
 OAI21_X2 _27879_ (.A(_04844_),
    .B1(_04846_),
    .B2(_04341_),
    .ZN(_04847_));
 NOR3_X1 _27880_ (.A1(_04454_),
    .A2(_04733_),
    .A3(_04479_),
    .ZN(_04848_));
 OR3_X1 _27881_ (.A1(_04521_),
    .A2(_04513_),
    .A3(_04848_),
    .ZN(_04849_));
 MUX2_X1 _27882_ (.A(net1198),
    .B(_04235_),
    .S(_04268_),
    .Z(_04850_));
 OAI221_X1 _27883_ (.A(_04460_),
    .B1(_04850_),
    .B2(_04564_),
    .C1(_04380_),
    .C2(_04440_),
    .ZN(_04851_));
 AND4_X1 _27884_ (.A1(_04379_),
    .A2(_04847_),
    .A3(_04849_),
    .A4(_04851_),
    .ZN(_04852_));
 OAI33_X1 _27885_ (.A1(_04818_),
    .A2(_04825_),
    .A3(_04831_),
    .B1(_04852_),
    .B2(_04841_),
    .B3(_04836_),
    .ZN(_00143_));
 INV_X1 _27886_ (.A(_06346_),
    .ZN(_04853_));
 NOR2_X1 _27887_ (.A1(_04853_),
    .A2(_09730_),
    .ZN(_04854_));
 NOR2_X1 _27888_ (.A1(_06346_),
    .A2(_09730_),
    .ZN(_04855_));
 XNOR2_X2 _27889_ (.A(_13179_),
    .B(_13224_),
    .ZN(_04856_));
 XNOR2_X2 _27890_ (.A(_10437_),
    .B(net584),
    .ZN(_04857_));
 XNOR2_X2 _27891_ (.A(_04856_),
    .B(_04857_),
    .ZN(_04858_));
 MUX2_X2 _27892_ (.A(_04854_),
    .B(_04855_),
    .S(_04858_),
    .Z(_04859_));
 OR3_X2 _27893_ (.A1(_06346_),
    .A2(_09856_),
    .A3(_00482_),
    .ZN(_04860_));
 NAND3_X2 _27894_ (.A1(_06346_),
    .A2(_00991_),
    .A3(_00482_),
    .ZN(_04861_));
 NAND2_X4 _27895_ (.A1(_04860_),
    .A2(_04861_),
    .ZN(_04862_));
 NOR2_X4 _27896_ (.A1(_04862_),
    .A2(_04859_),
    .ZN(_04863_));
 INV_X8 _27897_ (.A(_04863_),
    .ZN(_04864_));
 BUF_X16 _27898_ (.A(_04864_),
    .Z(_04865_));
 BUF_X16 _27899_ (.A(_04865_),
    .Z(_15264_));
 XNOR2_X1 _27900_ (.A(_10439_),
    .B(net574),
    .ZN(_04866_));
 XOR2_X2 _27901_ (.A(_10432_),
    .B(_10506_),
    .Z(_04867_));
 NAND3_X1 _27902_ (.A1(_06330_),
    .A2(_09100_),
    .A3(_04867_),
    .ZN(_04868_));
 NOR2_X1 _27903_ (.A1(_06330_),
    .A2(_08993_),
    .ZN(_04869_));
 NAND2_X1 _27904_ (.A1(_13224_),
    .A2(_04869_),
    .ZN(_04870_));
 AOI21_X1 _27905_ (.A(_04866_),
    .B1(_04868_),
    .B2(_04870_),
    .ZN(_04871_));
 XOR2_X1 _27906_ (.A(_10439_),
    .B(net573),
    .Z(_04872_));
 NAND2_X1 _27907_ (.A1(_04867_),
    .A2(_04869_),
    .ZN(_04873_));
 NAND3_X1 _27908_ (.A1(_06330_),
    .A2(_09023_),
    .A3(_13224_),
    .ZN(_04874_));
 AOI21_X1 _27909_ (.A(_04872_),
    .B1(_04873_),
    .B2(_04874_),
    .ZN(_04875_));
 INV_X1 _27910_ (.A(_06330_),
    .ZN(_04876_));
 NAND3_X1 _27911_ (.A1(_04876_),
    .A2(_09030_),
    .A3(_00483_),
    .ZN(_04877_));
 NAND2_X1 _27912_ (.A1(_06330_),
    .A2(_09030_),
    .ZN(_04878_));
 OAI21_X1 _27913_ (.A(_04877_),
    .B1(_04878_),
    .B2(_00483_),
    .ZN(_04879_));
 OR3_X4 _27914_ (.A1(_04871_),
    .A2(_04875_),
    .A3(_04879_),
    .ZN(_04880_));
 INV_X8 _27915_ (.A(_04880_),
    .ZN(_04881_));
 BUF_X4 clone13 (.A(_07376_),
    .Z(net13));
 BUF_X4 _27917_ (.A(_04881_),
    .Z(_15267_));
 XNOR2_X1 _27918_ (.A(_10550_),
    .B(_10482_),
    .ZN(_04883_));
 XOR2_X2 _27919_ (.A(net1068),
    .B(net586),
    .Z(_04884_));
 NAND3_X1 _27920_ (.A1(_06358_),
    .A2(_09194_),
    .A3(_04884_),
    .ZN(_04885_));
 NOR2_X1 _27921_ (.A1(_06358_),
    .A2(_09726_),
    .ZN(_04886_));
 NAND2_X1 _27922_ (.A1(_13167_),
    .A2(_04886_),
    .ZN(_04887_));
 AOI21_X2 _27923_ (.A(_04883_),
    .B1(_04885_),
    .B2(_04887_),
    .ZN(_04888_));
 XNOR2_X1 _27924_ (.A(_10550_),
    .B(_10480_),
    .ZN(_04889_));
 NAND2_X1 _27925_ (.A1(_04884_),
    .A2(_04886_),
    .ZN(_04890_));
 NAND3_X1 _27926_ (.A1(_06358_),
    .A2(_09074_),
    .A3(_13167_),
    .ZN(_04891_));
 AOI21_X2 _27927_ (.A(_04889_),
    .B1(_04890_),
    .B2(_04891_),
    .ZN(_04892_));
 NAND3_X1 _27928_ (.A1(_06365_),
    .A2(_08973_),
    .A3(_00484_),
    .ZN(_04893_));
 NAND2_X1 _27929_ (.A1(_06358_),
    .A2(_08973_),
    .ZN(_04894_));
 OAI21_X2 _27930_ (.A(_04893_),
    .B1(_04894_),
    .B2(_00484_),
    .ZN(_04895_));
 NOR3_X4 _27931_ (.A1(_04892_),
    .A2(_04888_),
    .A3(_04895_),
    .ZN(_04896_));
 INV_X4 _27932_ (.A(_04896_),
    .ZN(_04897_));
 BUF_X4 _27933_ (.A(_04897_),
    .Z(_04898_));
 BUF_X4 _27934_ (.A(_04898_),
    .Z(_04899_));
 BUF_X8 _27935_ (.A(_04899_),
    .Z(_04900_));
 BUF_X8 _27936_ (.A(_04900_),
    .Z(_15283_));
 BUF_X4 _27937_ (.A(_04880_),
    .Z(_04901_));
 BUF_X4 _27938_ (.A(_04901_),
    .Z(_15258_));
 BUF_X8 _27939_ (.A(_04896_),
    .Z(_04902_));
 BUF_X4 _27940_ (.A(_04902_),
    .Z(_04903_));
 BUF_X4 _27941_ (.A(_04903_),
    .Z(_04904_));
 BUF_X4 _27942_ (.A(_04904_),
    .Z(_04905_));
 BUF_X8 _27943_ (.A(_04905_),
    .Z(_15276_));
 XNOR2_X1 _27944_ (.A(_10503_),
    .B(_13229_),
    .ZN(_04906_));
 XNOR2_X2 _27945_ (.A(_10458_),
    .B(_04906_),
    .ZN(_04907_));
 MUX2_X2 _27946_ (.A(\text_in_r[39] ),
    .B(_04907_),
    .S(_11207_),
    .Z(_04908_));
 XOR2_X2 _27947_ (.A(_06442_),
    .B(_04908_),
    .Z(_04909_));
 XNOR2_X1 _27948_ (.A(_10516_),
    .B(_10505_),
    .ZN(_04910_));
 XNOR2_X2 _27949_ (.A(_10514_),
    .B(_04910_),
    .ZN(_04911_));
 XNOR2_X2 _27950_ (.A(_10524_),
    .B(_04911_),
    .ZN(_04912_));
 MUX2_X2 _27951_ (.A(\text_in_r[38] ),
    .B(_04912_),
    .S(_09803_),
    .Z(_04913_));
 XNOR2_X2 _27952_ (.A(_06434_),
    .B(_04913_),
    .ZN(_04914_));
 BUF_X4 _27953_ (.A(_04914_),
    .Z(_04915_));
 NOR2_X2 _27954_ (.A1(_04909_),
    .A2(_04915_),
    .ZN(_04916_));
 XNOR2_X1 _27955_ (.A(_10527_),
    .B(_10523_),
    .ZN(_04917_));
 XNOR2_X1 _27956_ (.A(_02320_),
    .B(_04917_),
    .ZN(_04918_));
 MUX2_X2 _27957_ (.A(\text_in_r[37] ),
    .B(_04918_),
    .S(_09076_),
    .Z(_04919_));
 XOR2_X2 _27958_ (.A(_06420_),
    .B(_04919_),
    .Z(_04920_));
 BUF_X4 _27959_ (.A(_04920_),
    .Z(_04921_));
 INV_X1 _27960_ (.A(_06406_),
    .ZN(_04922_));
 NOR2_X1 _27961_ (.A1(_09195_),
    .A2(\text_in_r[36] ),
    .ZN(_04923_));
 XNOR2_X1 _27962_ (.A(_10538_),
    .B(_02358_),
    .ZN(_04924_));
 AOI211_X2 _27963_ (.A(_04922_),
    .B(_04923_),
    .C1(_04924_),
    .C2(_11191_),
    .ZN(_04925_));
 AND2_X1 _27964_ (.A1(_11841_),
    .A2(\text_in_r[36] ),
    .ZN(_04926_));
 XOR2_X2 _27965_ (.A(_10538_),
    .B(_02358_),
    .Z(_04927_));
 AOI211_X2 _27966_ (.A(_06406_),
    .B(_04926_),
    .C1(_11191_),
    .C2(_04927_),
    .ZN(_04928_));
 OR2_X1 _27967_ (.A1(_04925_),
    .A2(_04928_),
    .ZN(_04929_));
 BUF_X2 _27968_ (.A(_04929_),
    .Z(_04930_));
 BUF_X4 _27969_ (.A(_04930_),
    .Z(_04931_));
 BUF_X4 _27970_ (.A(_04931_),
    .Z(_04932_));
 NAND2_X2 _27971_ (.A1(_04921_),
    .A2(_04932_),
    .ZN(_04933_));
 INV_X2 clone161 (.A(net10),
    .ZN(net161));
 BUF_X8 _27973_ (.A(net817),
    .Z(_04935_));
 AND2_X1 _27974_ (.A1(_06392_),
    .A2(net949),
    .ZN(_04936_));
 NOR2_X1 _27975_ (.A1(_06392_),
    .A2(_08994_),
    .ZN(_04937_));
 XNOR2_X2 _27976_ (.A(_10553_),
    .B(_02336_),
    .ZN(_04938_));
 MUX2_X1 _27977_ (.A(_04936_),
    .B(_04937_),
    .S(_04938_),
    .Z(_04939_));
 BUF_X8 _27978_ (.A(_04939_),
    .Z(_04940_));
 BUF_X2 _27979_ (.A(\text_in_r[35] ),
    .Z(_04941_));
 NOR2_X2 _27980_ (.A1(_06392_),
    .A2(_09075_),
    .ZN(_04942_));
 NAND2_X1 _27981_ (.A1(_04941_),
    .A2(_04942_),
    .ZN(_04943_));
 NAND2_X1 _27982_ (.A1(_06392_),
    .A2(_09730_),
    .ZN(_04944_));
 OAI21_X2 _27983_ (.A(_04943_),
    .B1(_04944_),
    .B2(_04941_),
    .ZN(_04945_));
 BUF_X8 _27984_ (.A(_04945_),
    .Z(_04946_));
 OAI21_X4 _27985_ (.A(_04896_),
    .B1(_04940_),
    .B2(_04946_),
    .ZN(_04947_));
 NAND2_X1 _27986_ (.A1(_04901_),
    .A2(_04897_),
    .ZN(_04948_));
 INV_X1 _27987_ (.A(_04936_),
    .ZN(_04949_));
 INV_X1 _27988_ (.A(_04937_),
    .ZN(_04950_));
 MUX2_X2 _27989_ (.A(_04949_),
    .B(_04950_),
    .S(_04938_),
    .Z(_04951_));
 BUF_X4 _27990_ (.A(_04951_),
    .Z(_04952_));
 NOR2_X1 _27991_ (.A1(_04941_),
    .A2(_04944_),
    .ZN(_04953_));
 AOI21_X4 _27992_ (.A(_04953_),
    .B1(_04942_),
    .B2(_04941_),
    .ZN(_04954_));
 BUF_X8 _27993_ (.A(_04954_),
    .Z(_04955_));
 AOI211_X2 _27994_ (.A(_04859_),
    .B(_04862_),
    .C1(_04952_),
    .C2(_04955_),
    .ZN(_04956_));
 OAI22_X1 _27995_ (.A1(net1113),
    .A2(_04947_),
    .B1(_04948_),
    .B2(_04956_),
    .ZN(_04957_));
 BUF_X8 _27996_ (.A(_04940_),
    .Z(_04958_));
 BUF_X8 _27997_ (.A(_04946_),
    .Z(_04959_));
 NOR3_X4 _27998_ (.A1(_04901_),
    .A2(_04958_),
    .A3(_04959_),
    .ZN(_04960_));
 NAND2_X1 _27999_ (.A1(_06346_),
    .A2(_09138_),
    .ZN(_04961_));
 NAND2_X1 _28000_ (.A1(_04853_),
    .A2(_09138_),
    .ZN(_04962_));
 MUX2_X2 _28001_ (.A(_04961_),
    .B(_04962_),
    .S(_04858_),
    .Z(_04963_));
 AND2_X1 _28002_ (.A1(_04860_),
    .A2(_04861_),
    .ZN(_04964_));
 NAND4_X2 _28003_ (.A1(_04963_),
    .A2(_04964_),
    .A3(_04951_),
    .A4(_04954_),
    .ZN(_04965_));
 BUF_X4 _28004_ (.A(_04965_),
    .Z(_04966_));
 CLKBUF_X2 split97 (.A(net709),
    .Z(net97));
 OAI21_X4 _28006_ (.A(net709),
    .B1(_04958_),
    .B2(_04959_),
    .ZN(_04968_));
 NAND2_X1 _28007_ (.A1(_04966_),
    .A2(_04968_),
    .ZN(_04969_));
 BUF_X4 _28008_ (.A(_04898_),
    .Z(_04970_));
 BUF_X4 _28009_ (.A(_04970_),
    .Z(_04971_));
 BUF_X4 _28010_ (.A(_15261_),
    .Z(_04972_));
 BUF_X8 _28011_ (.A(_04972_),
    .Z(_04973_));
 AOI21_X2 _28012_ (.A(_04897_),
    .B1(_04952_),
    .B2(_04955_),
    .ZN(_04974_));
 BUF_X4 _28013_ (.A(_04974_),
    .Z(_04975_));
 AOI221_X2 _28014_ (.A(_04960_),
    .B1(_04969_),
    .B2(_04971_),
    .C1(net1155),
    .C2(_04975_),
    .ZN(_04976_));
 NOR2_X4 _28015_ (.A1(_04925_),
    .A2(net1150),
    .ZN(_04977_));
 NAND2_X4 _28016_ (.A1(_04920_),
    .A2(_04977_),
    .ZN(_04978_));
 OAI221_X2 _28017_ (.A(_04916_),
    .B1(_04933_),
    .B2(_04957_),
    .C1(_04976_),
    .C2(_04978_),
    .ZN(_04979_));
 BUF_X4 _28018_ (.A(_04921_),
    .Z(_04980_));
 BUF_X4 _28019_ (.A(_04977_),
    .Z(_04981_));
 BUF_X4 _28020_ (.A(_04981_),
    .Z(_04982_));
 CLKBUF_X3 _28021_ (.A(_04970_),
    .Z(_04983_));
 NAND3_X1 _28022_ (.A1(_15258_),
    .A2(_04983_),
    .A3(_04966_),
    .ZN(_04984_));
 NAND2_X4 _28023_ (.A1(_04952_),
    .A2(_04955_),
    .ZN(_04985_));
 CLKBUF_X3 _28024_ (.A(_04985_),
    .Z(_04986_));
 BUF_X16 _28025_ (.A(_04863_),
    .Z(_04987_));
 BUF_X4 clone650 (.A(net817),
    .Z(net1113));
 OAI21_X1 _28027_ (.A(_04968_),
    .B1(_04986_),
    .B2(net95),
    .ZN(_04989_));
 OAI21_X1 _28028_ (.A(_04984_),
    .B1(_04989_),
    .B2(_04971_),
    .ZN(_04990_));
 CLKBUF_X3 _28029_ (.A(_04930_),
    .Z(_04991_));
 BUF_X4 _28030_ (.A(_04991_),
    .Z(_04992_));
 NAND2_X4 _28031_ (.A1(_04881_),
    .A2(_04896_),
    .ZN(_04993_));
 OAI221_X2 _28032_ (.A(_04948_),
    .B1(_04993_),
    .B2(_04987_),
    .C1(_04958_),
    .C2(_04959_),
    .ZN(_04994_));
 AND2_X1 _28033_ (.A1(_04992_),
    .A2(_04994_),
    .ZN(_04995_));
 OAI21_X4 _28034_ (.A(_04970_),
    .B1(_04862_),
    .B2(net507),
    .ZN(_04996_));
 BUF_X4 _28035_ (.A(_04985_),
    .Z(_04997_));
 BUF_X4 _28036_ (.A(_04997_),
    .Z(_04998_));
 BUF_X1 split32 (.A(_14694_),
    .Z(net32));
 INV_X1 _28038_ (.A(net896),
    .ZN(_05000_));
 AOI21_X1 _28039_ (.A(_04998_),
    .B1(_04905_),
    .B2(_05000_),
    .ZN(_05001_));
 NAND2_X1 _28040_ (.A1(_04996_),
    .A2(_05001_),
    .ZN(_05002_));
 AOI221_X2 _28041_ (.A(_04980_),
    .B1(_04982_),
    .B2(_04990_),
    .C1(_04995_),
    .C2(_05002_),
    .ZN(_05003_));
 BUF_X4 _28042_ (.A(_04909_),
    .Z(_05004_));
 XOR2_X2 _28043_ (.A(_06434_),
    .B(_04913_),
    .Z(_05005_));
 NAND2_X2 _28044_ (.A1(_05004_),
    .A2(_05005_),
    .ZN(_05006_));
 BUF_X2 _28045_ (.A(_15260_),
    .Z(_05007_));
 CLKBUF_X3 _28046_ (.A(_05007_),
    .Z(_05008_));
 INV_X1 _28047_ (.A(_05008_),
    .ZN(_05009_));
 NAND3_X1 _28048_ (.A1(_04897_),
    .A2(_04951_),
    .A3(_04954_),
    .ZN(_05010_));
 CLKBUF_X3 _28049_ (.A(_05010_),
    .Z(_05011_));
 OR2_X1 _28050_ (.A1(_05009_),
    .A2(_05011_),
    .ZN(_05012_));
 AOI21_X4 _28051_ (.A(net817),
    .B1(_04952_),
    .B2(_04955_),
    .ZN(_05013_));
 NOR3_X4 _28052_ (.A1(net896),
    .A2(_04940_),
    .A3(_04946_),
    .ZN(_05014_));
 OAI21_X1 _28053_ (.A(_04903_),
    .B1(_05013_),
    .B2(_05014_),
    .ZN(_05015_));
 AOI21_X2 _28054_ (.A(_04978_),
    .B1(_05012_),
    .B2(_05015_),
    .ZN(_05016_));
 NOR2_X4 _28055_ (.A1(_04940_),
    .A2(_04946_),
    .ZN(_05017_));
 BUF_X4 _28056_ (.A(_05017_),
    .Z(_05018_));
 BUF_X4 _28057_ (.A(_05018_),
    .Z(_05019_));
 AND2_X2 _28058_ (.A1(net818),
    .A2(_04898_),
    .ZN(_05020_));
 AOI21_X1 _28059_ (.A(_04921_),
    .B1(_05019_),
    .B2(_05020_),
    .ZN(_05021_));
 BUF_X4 clone6 (.A(_06216_),
    .Z(net6));
 INV_X4 _28061_ (.A(_15270_),
    .ZN(_05023_));
 NOR2_X1 _28062_ (.A1(_05023_),
    .A2(_04898_),
    .ZN(_05024_));
 OAI22_X1 _28063_ (.A1(_04973_),
    .A2(_04947_),
    .B1(_05024_),
    .B2(_04997_),
    .ZN(_05025_));
 MUX2_X1 _28064_ (.A(_04994_),
    .B(_05025_),
    .S(_04981_),
    .Z(_05026_));
 NAND2_X4 _28065_ (.A1(net698),
    .A2(_04898_),
    .ZN(_05027_));
 OAI21_X4 _28066_ (.A(_04902_),
    .B1(_04862_),
    .B2(_04859_),
    .ZN(_05028_));
 NAND3_X1 _28067_ (.A1(_05018_),
    .A2(_05027_),
    .A3(_05028_),
    .ZN(_05029_));
 NOR2_X4 _28068_ (.A1(_04880_),
    .A2(_04897_),
    .ZN(_05030_));
 BUF_X4 clone159 (.A(_04864_),
    .Z(net159));
 NOR2_X1 _28070_ (.A1(net160),
    .A2(_04903_),
    .ZN(_05032_));
 OAI21_X1 _28071_ (.A(_04986_),
    .B1(_05030_),
    .B2(_05032_),
    .ZN(_05033_));
 AND3_X1 _28072_ (.A1(_04932_),
    .A2(_05029_),
    .A3(_05033_),
    .ZN(_05034_));
 AOI221_X2 _28073_ (.A(_05016_),
    .B1(_05026_),
    .B2(_05021_),
    .C1(_04980_),
    .C2(_05034_),
    .ZN(_05035_));
 OAI22_X2 _28074_ (.A1(_04979_),
    .A2(_05003_),
    .B1(_05035_),
    .B2(_05006_),
    .ZN(_05036_));
 NAND2_X2 _28075_ (.A1(_05004_),
    .A2(_04915_),
    .ZN(_05037_));
 BUF_X4 _28076_ (.A(_04981_),
    .Z(_05038_));
 BUF_X4 _28077_ (.A(_04865_),
    .Z(_05039_));
 NOR2_X4 _28078_ (.A1(_04881_),
    .A2(net1148),
    .ZN(_05040_));
 BUF_X4 _28079_ (.A(_04952_),
    .Z(_05041_));
 BUF_X8 _28080_ (.A(_04955_),
    .Z(_05042_));
 NAND3_X4 _28081_ (.A1(net817),
    .A2(_05041_),
    .A3(_05042_),
    .ZN(_05043_));
 NAND3_X4 _28082_ (.A1(_04896_),
    .A2(_04951_),
    .A3(_04954_),
    .ZN(_05044_));
 AOI22_X2 _28083_ (.A1(_05039_),
    .A2(_05040_),
    .B1(_05043_),
    .B2(_05044_),
    .ZN(_05045_));
 NOR2_X2 _28084_ (.A1(_05007_),
    .A2(_04947_),
    .ZN(_05046_));
 NOR3_X2 _28085_ (.A1(_05038_),
    .A2(_05045_),
    .A3(_05046_),
    .ZN(_05047_));
 NAND3_X2 _28086_ (.A1(net897),
    .A2(_05041_),
    .A3(_05042_),
    .ZN(_05048_));
 OAI21_X4 _28087_ (.A(_04881_),
    .B1(_04958_),
    .B2(_04959_),
    .ZN(_05049_));
 AND2_X1 _28088_ (.A1(_05048_),
    .A2(_05049_),
    .ZN(_05050_));
 BUF_X4 _28089_ (.A(_04904_),
    .Z(_05051_));
 OAI21_X1 _28090_ (.A(_05047_),
    .B1(_05050_),
    .B2(_05051_),
    .ZN(_05052_));
 NOR2_X1 _28091_ (.A1(_04903_),
    .A2(_04985_),
    .ZN(_05053_));
 AOI221_X2 _28092_ (.A(_04931_),
    .B1(_04997_),
    .B2(_15281_),
    .C1(_05053_),
    .C2(net1155),
    .ZN(_05054_));
 NOR2_X1 _28093_ (.A1(_04980_),
    .A2(_05054_),
    .ZN(_05055_));
 BUF_X4 _28094_ (.A(_04932_),
    .Z(_05056_));
 NAND2_X2 _28095_ (.A1(_04901_),
    .A2(_04902_),
    .ZN(_05057_));
 NOR2_X2 _28096_ (.A1(net94),
    .A2(_05057_),
    .ZN(_05058_));
 OAI21_X4 _28097_ (.A(_15270_),
    .B1(_04958_),
    .B2(_04959_),
    .ZN(_05059_));
 MUX2_X1 _28098_ (.A(_05000_),
    .B(_05058_),
    .S(_04986_),
    .Z(_05060_));
 CLKBUF_X3 _28099_ (.A(_04983_),
    .Z(_05061_));
 OAI221_X2 _28100_ (.A(_05056_),
    .B1(_05058_),
    .B2(_05059_),
    .C1(_05060_),
    .C2(_05061_),
    .ZN(_05062_));
 XNOR2_X2 _28101_ (.A(_06420_),
    .B(_04919_),
    .ZN(_05063_));
 BUF_X4 _28102_ (.A(_05063_),
    .Z(_05064_));
 BUF_X4 _28103_ (.A(_05064_),
    .Z(_05065_));
 AOI21_X1 _28104_ (.A(_04986_),
    .B1(_05040_),
    .B2(_05039_),
    .ZN(_05066_));
 BUF_X4 _28105_ (.A(_05017_),
    .Z(_05067_));
 BUF_X4 _28106_ (.A(_05067_),
    .Z(_05068_));
 NOR2_X1 _28107_ (.A1(_05000_),
    .A2(_05068_),
    .ZN(_05069_));
 OAI21_X1 _28108_ (.A(_05051_),
    .B1(_05066_),
    .B2(_05069_),
    .ZN(_05070_));
 INV_X2 _28109_ (.A(_15268_),
    .ZN(_05071_));
 AOI21_X1 _28110_ (.A(_04992_),
    .B1(_05066_),
    .B2(_05071_),
    .ZN(_05072_));
 AOI21_X1 _28111_ (.A(_05065_),
    .B1(_05070_),
    .B2(_05072_),
    .ZN(_05073_));
 AOI221_X2 _28112_ (.A(_05037_),
    .B1(_05052_),
    .B2(_05055_),
    .C1(_05062_),
    .C2(_05073_),
    .ZN(_05074_));
 BUF_X4 _28113_ (.A(_04980_),
    .Z(_05075_));
 AOI21_X2 _28114_ (.A(_04997_),
    .B1(_04881_),
    .B2(_04865_),
    .ZN(_05076_));
 OAI21_X1 _28115_ (.A(_05061_),
    .B1(_05019_),
    .B2(_05008_),
    .ZN(_05077_));
 NAND3_X4 _28116_ (.A1(_04972_),
    .A2(_04952_),
    .A3(_04955_),
    .ZN(_05078_));
 BUF_X4 _28117_ (.A(_05019_),
    .Z(_05079_));
 OAI21_X1 _28118_ (.A(_05078_),
    .B1(_05079_),
    .B2(net160),
    .ZN(_05080_));
 OAI221_X1 _28119_ (.A(_05075_),
    .B1(_05076_),
    .B2(_05077_),
    .C1(_05080_),
    .C2(_15283_),
    .ZN(_05081_));
 NOR2_X1 _28120_ (.A1(net160),
    .A2(_05011_),
    .ZN(_05082_));
 OAI21_X4 _28121_ (.A(net1148),
    .B1(_04958_),
    .B2(_04959_),
    .ZN(_05083_));
 NAND2_X1 _28122_ (.A1(_05044_),
    .A2(_05083_),
    .ZN(_05084_));
 AOI221_X1 _28123_ (.A(_05082_),
    .B1(_05084_),
    .B2(_05009_),
    .C1(_04975_),
    .C2(net1155),
    .ZN(_05085_));
 OAI21_X1 _28124_ (.A(_05081_),
    .B1(_05085_),
    .B2(_05075_),
    .ZN(_05086_));
 BUF_X4 _28125_ (.A(_04992_),
    .Z(_05087_));
 NOR2_X1 _28126_ (.A1(_05004_),
    .A2(_05005_),
    .ZN(_05088_));
 NAND2_X1 _28127_ (.A1(_05087_),
    .A2(_05088_),
    .ZN(_05089_));
 NAND2_X1 _28128_ (.A1(_04982_),
    .A2(_05088_),
    .ZN(_05090_));
 NOR2_X1 _28129_ (.A1(_04904_),
    .A2(_04920_),
    .ZN(_05091_));
 INV_X8 _28130_ (.A(_04972_),
    .ZN(_05092_));
 OAI21_X1 _28131_ (.A(_04993_),
    .B1(_04881_),
    .B2(_05039_),
    .ZN(_05093_));
 AOI221_X1 _28132_ (.A(_05068_),
    .B1(_05091_),
    .B2(net1157),
    .C1(_05093_),
    .C2(_04921_),
    .ZN(_05094_));
 NOR3_X1 _28133_ (.A1(net1157),
    .A2(_04899_),
    .A3(_04920_),
    .ZN(_05095_));
 NOR2_X4 _28134_ (.A1(_04880_),
    .A2(_04896_),
    .ZN(_05096_));
 OAI21_X1 _28135_ (.A(_04904_),
    .B1(_05064_),
    .B2(_04881_),
    .ZN(_05097_));
 AOI221_X2 _28136_ (.A(_05095_),
    .B1(_05096_),
    .B2(_04921_),
    .C1(_15264_),
    .C2(_05097_),
    .ZN(_05098_));
 AOI21_X1 _28137_ (.A(_05094_),
    .B1(_05098_),
    .B2(_05079_),
    .ZN(_05099_));
 OAI22_X2 _28138_ (.A1(_05086_),
    .A2(_05089_),
    .B1(_05090_),
    .B2(_05099_),
    .ZN(_05100_));
 NOR3_X4 _28139_ (.A1(_05036_),
    .A2(_05074_),
    .A3(_05100_),
    .ZN(_00144_));
 BUF_X4 _28140_ (.A(_05063_),
    .Z(_05101_));
 NAND2_X1 _28141_ (.A1(_05039_),
    .A2(_04960_),
    .ZN(_05102_));
 AOI22_X1 _28142_ (.A1(_04983_),
    .A2(_04968_),
    .B1(_04975_),
    .B2(net95),
    .ZN(_05103_));
 NAND3_X1 _28143_ (.A1(_04982_),
    .A2(_05102_),
    .A3(_05103_),
    .ZN(_05104_));
 BUF_X4 _28144_ (.A(_04903_),
    .Z(_05105_));
 OAI21_X4 _28145_ (.A(_05092_),
    .B1(_04940_),
    .B2(_04946_),
    .ZN(_05106_));
 NAND3_X1 _28146_ (.A1(_05105_),
    .A2(_05043_),
    .A3(net1112),
    .ZN(_05107_));
 AOI21_X2 _28147_ (.A(_05017_),
    .B1(_04881_),
    .B2(_04865_),
    .ZN(_05108_));
 OAI221_X2 _28148_ (.A(_05107_),
    .B1(net1151),
    .B2(_04925_),
    .C1(_04905_),
    .C2(_05108_),
    .ZN(_05109_));
 AOI21_X1 _28149_ (.A(_05101_),
    .B1(_05104_),
    .B2(_05109_),
    .ZN(_05110_));
 NOR2_X2 _28150_ (.A1(_04920_),
    .A2(_04977_),
    .ZN(_05111_));
 OAI221_X1 _28151_ (.A(_05111_),
    .B1(_05049_),
    .B2(_05039_),
    .C1(net1157),
    .C2(_05011_),
    .ZN(_05112_));
 AOI21_X1 _28152_ (.A(_05112_),
    .B1(_05084_),
    .B2(_15258_),
    .ZN(_05113_));
 NAND2_X2 _28153_ (.A1(_05064_),
    .A2(_04981_),
    .ZN(_05114_));
 OAI21_X4 _28154_ (.A(_04972_),
    .B1(_04940_),
    .B2(_04946_),
    .ZN(_05115_));
 NAND3_X4 _28155_ (.A1(_05007_),
    .A2(_05041_),
    .A3(_05042_),
    .ZN(_05116_));
 AOI21_X1 _28156_ (.A(_04983_),
    .B1(_05115_),
    .B2(_05116_),
    .ZN(_05117_));
 AOI21_X1 _28157_ (.A(_04960_),
    .B1(_04997_),
    .B2(net818),
    .ZN(_05118_));
 AND2_X1 _28158_ (.A1(_04983_),
    .A2(_05118_),
    .ZN(_05119_));
 NOR3_X1 _28159_ (.A1(_05114_),
    .A2(_05117_),
    .A3(_05119_),
    .ZN(_05120_));
 NOR4_X2 _28160_ (.A1(_05006_),
    .A2(_05110_),
    .A3(_05113_),
    .A4(_05120_),
    .ZN(_05121_));
 AOI21_X1 _28161_ (.A(_04900_),
    .B1(net1112),
    .B2(_05102_),
    .ZN(_05122_));
 OAI21_X1 _28162_ (.A(_05111_),
    .B1(_05011_),
    .B2(_15267_),
    .ZN(_05123_));
 OAI21_X1 _28163_ (.A(_04916_),
    .B1(_05122_),
    .B2(_05123_),
    .ZN(_05124_));
 NOR3_X1 _28164_ (.A1(_04987_),
    .A2(_04901_),
    .A3(_05067_),
    .ZN(_05125_));
 OR3_X1 _28165_ (.A1(_04905_),
    .A2(_05014_),
    .A3(_05125_),
    .ZN(_05126_));
 CLKBUF_X3 _28166_ (.A(_04998_),
    .Z(_05127_));
 OAI21_X1 _28167_ (.A(_05115_),
    .B1(_05127_),
    .B2(net97),
    .ZN(_05128_));
 OAI21_X1 _28168_ (.A(_05126_),
    .B1(_05128_),
    .B2(_05061_),
    .ZN(_05129_));
 NOR2_X1 _28169_ (.A1(_04980_),
    .A2(_05056_),
    .ZN(_05130_));
 AOI21_X1 _28170_ (.A(_05124_),
    .B1(_05129_),
    .B2(_05130_),
    .ZN(_05131_));
 NAND3_X4 _28171_ (.A1(_04881_),
    .A2(_05041_),
    .A3(_05042_),
    .ZN(_05132_));
 AOI21_X2 _28172_ (.A(_04904_),
    .B1(_05132_),
    .B2(_05115_),
    .ZN(_05133_));
 AOI21_X1 _28173_ (.A(_05014_),
    .B1(_04998_),
    .B2(_05008_),
    .ZN(_05134_));
 AOI21_X1 _28174_ (.A(_05133_),
    .B1(_05134_),
    .B2(_05051_),
    .ZN(_05135_));
 NOR2_X1 _28175_ (.A1(_05056_),
    .A2(_05135_),
    .ZN(_05136_));
 OAI21_X1 _28176_ (.A(_05105_),
    .B1(_04960_),
    .B2(net816),
    .ZN(_05137_));
 OAI21_X1 _28177_ (.A(_05116_),
    .B1(_05068_),
    .B2(_05039_),
    .ZN(_05138_));
 NAND2_X1 _28178_ (.A1(_04900_),
    .A2(_05138_),
    .ZN(_05139_));
 AND3_X1 _28179_ (.A1(_04992_),
    .A2(_05137_),
    .A3(_05139_),
    .ZN(_05140_));
 OAI21_X1 _28180_ (.A(_05075_),
    .B1(_05136_),
    .B2(_05140_),
    .ZN(_05141_));
 XNOR2_X2 _28181_ (.A(_06442_),
    .B(_04908_),
    .ZN(_05142_));
 BUF_X4 _28182_ (.A(_05142_),
    .Z(_05143_));
 AOI221_X2 _28183_ (.A(_04985_),
    .B1(_05030_),
    .B2(_04864_),
    .C1(_04898_),
    .C2(_15268_),
    .ZN(_05144_));
 NAND2_X1 _28184_ (.A1(_05008_),
    .A2(_04970_),
    .ZN(_05145_));
 AOI21_X1 _28185_ (.A(_04986_),
    .B1(_05057_),
    .B2(_05145_),
    .ZN(_05146_));
 NOR2_X1 _28186_ (.A1(_05040_),
    .A2(_05096_),
    .ZN(_05147_));
 NOR2_X1 _28187_ (.A1(net95),
    .A2(_05018_),
    .ZN(_05148_));
 AOI21_X1 _28188_ (.A(_05146_),
    .B1(_05147_),
    .B2(_05148_),
    .ZN(_05149_));
 MUX2_X1 _28189_ (.A(_05144_),
    .B(_05149_),
    .S(_05038_),
    .Z(_05150_));
 NOR2_X1 _28190_ (.A1(_15284_),
    .A2(_05068_),
    .ZN(_05151_));
 NOR3_X1 _28191_ (.A1(_04982_),
    .A2(_05144_),
    .A3(_05151_),
    .ZN(_05152_));
 NOR2_X1 _28192_ (.A1(_04980_),
    .A2(_05152_),
    .ZN(_05153_));
 AOI211_X2 _28193_ (.A(_04940_),
    .B(_04946_),
    .C1(_04963_),
    .C2(_04964_),
    .ZN(_05154_));
 OAI21_X1 _28194_ (.A(_04900_),
    .B1(_05154_),
    .B2(_04956_),
    .ZN(_05155_));
 AND2_X1 _28195_ (.A1(_05155_),
    .A2(_05137_),
    .ZN(_05156_));
 OAI221_X2 _28196_ (.A(_05143_),
    .B1(_05150_),
    .B2(_05153_),
    .C1(_05114_),
    .C2(_05156_),
    .ZN(_05157_));
 NAND3_X1 _28197_ (.A1(_04977_),
    .A2(_05067_),
    .A3(_05096_),
    .ZN(_05158_));
 NAND3_X1 _28198_ (.A1(_04920_),
    .A2(_04909_),
    .A3(_05158_),
    .ZN(_05159_));
 NAND2_X2 _28199_ (.A1(_04977_),
    .A2(_05067_),
    .ZN(_05160_));
 NOR2_X1 _28200_ (.A1(_05092_),
    .A2(_04930_),
    .ZN(_05161_));
 OAI22_X1 _28201_ (.A1(_04935_),
    .A2(_05160_),
    .B1(_05161_),
    .B2(_05018_),
    .ZN(_05162_));
 AOI21_X2 _28202_ (.A(_05159_),
    .B1(_05162_),
    .B2(_05105_),
    .ZN(_05163_));
 NAND2_X1 _28203_ (.A1(_04898_),
    .A2(_04977_),
    .ZN(_05164_));
 OAI22_X2 _28204_ (.A1(_04981_),
    .A2(_04966_),
    .B1(_05164_),
    .B2(_05067_),
    .ZN(_05165_));
 OAI22_X1 _28205_ (.A1(_04899_),
    .A2(_04977_),
    .B1(_05083_),
    .B2(_04881_),
    .ZN(_05166_));
 AOI22_X2 _28206_ (.A1(_15258_),
    .A2(_05165_),
    .B1(_05166_),
    .B2(_05039_),
    .ZN(_05167_));
 AND2_X1 _28207_ (.A1(_05044_),
    .A2(_05083_),
    .ZN(_05168_));
 OAI221_X1 _28208_ (.A(_04981_),
    .B1(_05011_),
    .B2(_04935_),
    .C1(_05168_),
    .C2(net95),
    .ZN(_05169_));
 NAND3_X1 _28209_ (.A1(_04899_),
    .A2(_05043_),
    .A3(_05115_),
    .ZN(_05170_));
 NAND2_X2 _28210_ (.A1(net159),
    .A2(_05040_),
    .ZN(_05171_));
 OAI221_X1 _28211_ (.A(_05170_),
    .B1(_05171_),
    .B2(_04986_),
    .C1(net97),
    .C2(_04947_),
    .ZN(_05172_));
 OAI21_X1 _28212_ (.A(_05169_),
    .B1(_05172_),
    .B2(_05038_),
    .ZN(_05173_));
 NOR2_X1 _28213_ (.A1(_04980_),
    .A2(_05143_),
    .ZN(_05174_));
 AOI221_X2 _28214_ (.A(_05005_),
    .B1(_05163_),
    .B2(_05167_),
    .C1(_05173_),
    .C2(_05174_),
    .ZN(_05175_));
 AOI221_X2 _28215_ (.A(_05121_),
    .B1(_05141_),
    .B2(_05131_),
    .C1(_05157_),
    .C2(_05175_),
    .ZN(_00145_));
 NOR2_X1 _28216_ (.A1(_05101_),
    .A2(_05056_),
    .ZN(_05176_));
 NOR3_X4 _28217_ (.A1(_15274_),
    .A2(_04940_),
    .A3(_04946_),
    .ZN(_05177_));
 OAI21_X1 _28218_ (.A(_15283_),
    .B1(_05148_),
    .B2(_05177_),
    .ZN(_05178_));
 NAND3_X1 _28219_ (.A1(_15276_),
    .A2(_05132_),
    .A3(_05059_),
    .ZN(_05179_));
 AND3_X1 _28220_ (.A1(_05176_),
    .A2(_05178_),
    .A3(_05179_),
    .ZN(_05180_));
 OR2_X1 _28221_ (.A1(_04935_),
    .A2(_05105_),
    .ZN(_05181_));
 NAND2_X1 _28222_ (.A1(_05111_),
    .A2(_05181_),
    .ZN(_05182_));
 NAND3_X2 _28223_ (.A1(net898),
    .A2(_05041_),
    .A3(_05042_),
    .ZN(_05183_));
 BUF_X32 _28224_ (.A(_04987_),
    .Z(_15259_));
 OAI21_X1 _28225_ (.A(_05183_),
    .B1(_05079_),
    .B2(net96),
    .ZN(_05184_));
 NOR2_X1 _28226_ (.A1(_15283_),
    .A2(_05184_),
    .ZN(_05185_));
 OAI21_X1 _28227_ (.A(_04916_),
    .B1(_05182_),
    .B2(_05185_),
    .ZN(_05186_));
 NOR2_X2 _28228_ (.A1(_05101_),
    .A2(_05038_),
    .ZN(_05187_));
 NAND3_X1 _28229_ (.A1(_15283_),
    .A2(net1112),
    .A3(_05183_),
    .ZN(_05188_));
 NAND3_X1 _28230_ (.A1(_15276_),
    .A2(_05132_),
    .A3(_05115_),
    .ZN(_05189_));
 NAND3_X1 _28231_ (.A1(_05187_),
    .A2(_05188_),
    .A3(_05189_),
    .ZN(_05190_));
 AOI21_X4 _28232_ (.A(_04881_),
    .B1(_04952_),
    .B2(_04955_),
    .ZN(_05191_));
 NOR3_X2 _28233_ (.A1(net188),
    .A2(_04958_),
    .A3(_04959_),
    .ZN(_05192_));
 NOR3_X1 _28234_ (.A1(_05061_),
    .A2(_05191_),
    .A3(_05192_),
    .ZN(_05193_));
 NOR3_X1 _28235_ (.A1(_15276_),
    .A2(net816),
    .A3(_05177_),
    .ZN(_05194_));
 OAI21_X1 _28236_ (.A(_05130_),
    .B1(_05193_),
    .B2(_05194_),
    .ZN(_05195_));
 NAND2_X1 _28237_ (.A1(_05190_),
    .A2(_05195_),
    .ZN(_05196_));
 NOR3_X1 _28238_ (.A1(_05180_),
    .A2(_05186_),
    .A3(_05196_),
    .ZN(_05197_));
 NAND2_X2 _28239_ (.A1(_05142_),
    .A2(_04915_),
    .ZN(_05198_));
 NOR2_X2 _28240_ (.A1(_04898_),
    .A2(_04985_),
    .ZN(_05199_));
 NAND3_X2 _28241_ (.A1(_15274_),
    .A2(_04952_),
    .A3(_04955_),
    .ZN(_05200_));
 NAND2_X1 _28242_ (.A1(_05049_),
    .A2(_05200_),
    .ZN(_05201_));
 AOI221_X2 _28243_ (.A(_04956_),
    .B1(_05199_),
    .B2(net1113),
    .C1(_05201_),
    .C2(_04971_),
    .ZN(_05202_));
 AOI21_X2 _28244_ (.A(_05079_),
    .B1(_05171_),
    .B2(_05181_),
    .ZN(_05203_));
 NAND2_X1 _28245_ (.A1(_05087_),
    .A2(_05029_),
    .ZN(_05204_));
 OAI221_X1 _28246_ (.A(_05065_),
    .B1(_05087_),
    .B2(_05202_),
    .C1(_05203_),
    .C2(_05204_),
    .ZN(_05205_));
 AOI21_X1 _28247_ (.A(_05061_),
    .B1(_05049_),
    .B2(_05078_),
    .ZN(_05206_));
 AOI21_X1 _28248_ (.A(net189),
    .B1(_05041_),
    .B2(_05042_),
    .ZN(_05207_));
 NOR3_X1 _28249_ (.A1(_05051_),
    .A2(_05154_),
    .A3(_05207_),
    .ZN(_05208_));
 NOR3_X1 _28250_ (.A1(_04978_),
    .A2(_05206_),
    .A3(_05208_),
    .ZN(_05209_));
 OAI33_X1 _28251_ (.A1(net97),
    .A2(_15283_),
    .A3(_05079_),
    .B1(_04960_),
    .B2(_04996_),
    .B3(_05191_),
    .ZN(_05210_));
 AOI21_X2 _28252_ (.A(_05209_),
    .B1(_05210_),
    .B2(_05187_),
    .ZN(_05211_));
 AOI21_X1 _28253_ (.A(_05198_),
    .B1(_05205_),
    .B2(_05211_),
    .ZN(_05212_));
 NOR3_X1 _28254_ (.A1(_15259_),
    .A2(_04932_),
    .A3(_05096_),
    .ZN(_05213_));
 AND2_X1 _28255_ (.A1(_15279_),
    .A2(_04991_),
    .ZN(_05214_));
 INV_X1 _28256_ (.A(_15288_),
    .ZN(_05215_));
 MUX2_X1 _28257_ (.A(_05215_),
    .B(_04986_),
    .S(_04931_),
    .Z(_05216_));
 OAI21_X2 _28258_ (.A(_04897_),
    .B1(_04925_),
    .B2(net1149),
    .ZN(_05217_));
 AOI221_X2 _28259_ (.A(_04881_),
    .B1(_05017_),
    .B2(_05217_),
    .C1(_04964_),
    .C2(_04963_),
    .ZN(_05218_));
 NOR2_X1 _28260_ (.A1(net1153),
    .A2(_04947_),
    .ZN(_05219_));
 OAI33_X1 _28261_ (.A1(_05079_),
    .A2(_05213_),
    .A3(_05214_),
    .B1(_05219_),
    .B2(_05218_),
    .B3(_05216_),
    .ZN(_05220_));
 AND2_X1 _28262_ (.A1(_05065_),
    .A2(_05220_),
    .ZN(_05221_));
 NOR2_X4 _28263_ (.A1(_15262_),
    .A2(net1114),
    .ZN(_05222_));
 OAI21_X1 _28264_ (.A(_04903_),
    .B1(_05067_),
    .B2(_05222_),
    .ZN(_05223_));
 NAND3_X2 _28265_ (.A1(_05071_),
    .A2(_05041_),
    .A3(_05042_),
    .ZN(_05224_));
 NAND2_X1 _28266_ (.A1(_04970_),
    .A2(_05224_),
    .ZN(_05225_));
 OAI22_X2 _28267_ (.A1(_05076_),
    .A2(_05223_),
    .B1(_05225_),
    .B2(_05108_),
    .ZN(_05226_));
 NAND3_X1 _28268_ (.A1(_04905_),
    .A2(net1112),
    .A3(_05116_),
    .ZN(_05227_));
 NOR2_X2 _28269_ (.A1(_04903_),
    .A2(_05017_),
    .ZN(_05228_));
 AOI21_X1 _28270_ (.A(_04981_),
    .B1(_05228_),
    .B2(net1113),
    .ZN(_05229_));
 AOI221_X2 _28271_ (.A(_05101_),
    .B1(_05038_),
    .B2(_05226_),
    .C1(_05227_),
    .C2(_05229_),
    .ZN(_05230_));
 OAI21_X2 _28272_ (.A(_15268_),
    .B1(_04958_),
    .B2(_04959_),
    .ZN(_05231_));
 NAND3_X1 _28273_ (.A1(_04905_),
    .A2(_04966_),
    .A3(_05231_),
    .ZN(_05232_));
 NAND3_X2 _28274_ (.A1(_05106_),
    .A2(_04971_),
    .A3(_05116_),
    .ZN(_05233_));
 AND3_X2 _28275_ (.A1(_05101_),
    .A2(_05232_),
    .A3(_05233_),
    .ZN(_05234_));
 NOR3_X1 _28276_ (.A1(net1153),
    .A2(_05068_),
    .A3(_05040_),
    .ZN(_05235_));
 NOR3_X1 _28277_ (.A1(_05039_),
    .A2(_04899_),
    .A3(_05191_),
    .ZN(_05236_));
 AOI21_X1 _28278_ (.A(_04973_),
    .B1(_04966_),
    .B2(_04996_),
    .ZN(_05237_));
 NOR4_X2 _28279_ (.A1(_05237_),
    .A2(_05235_),
    .A3(_05236_),
    .A4(_05101_),
    .ZN(_05238_));
 NOR3_X2 _28280_ (.A1(_05087_),
    .A2(_05234_),
    .A3(_05238_),
    .ZN(_05239_));
 OAI221_X2 _28281_ (.A(_05028_),
    .B1(_04959_),
    .B2(_04958_),
    .C1(_05039_),
    .C2(_04881_),
    .ZN(_05240_));
 INV_X1 _28282_ (.A(_15284_),
    .ZN(_05241_));
 AOI21_X1 _28283_ (.A(_04920_),
    .B1(_05018_),
    .B2(_05241_),
    .ZN(_05242_));
 NOR2_X2 _28284_ (.A1(net1156),
    .A2(_04902_),
    .ZN(_05243_));
 NOR2_X1 _28285_ (.A1(_05018_),
    .A2(_05243_),
    .ZN(_05244_));
 AOI22_X2 _28286_ (.A1(_15281_),
    .A2(_05068_),
    .B1(_05171_),
    .B2(_05244_),
    .ZN(_05245_));
 AOI221_X2 _28287_ (.A(_05038_),
    .B1(_05240_),
    .B2(_05242_),
    .C1(_05245_),
    .C2(_04921_),
    .ZN(_05246_));
 OAI33_X1 _28288_ (.A1(_05037_),
    .A2(_05221_),
    .A3(_05230_),
    .B1(_05006_),
    .B2(_05246_),
    .B3(_05239_),
    .ZN(_05247_));
 NOR3_X1 _28289_ (.A1(_05247_),
    .A2(_05212_),
    .A3(_05197_),
    .ZN(_00146_));
 NAND2_X1 _28290_ (.A1(_04902_),
    .A2(_04977_),
    .ZN(_05248_));
 MUX2_X1 _28291_ (.A(net1158),
    .B(_05092_),
    .S(_05217_),
    .Z(_05249_));
 NAND2_X1 _28292_ (.A1(_05248_),
    .A2(_05249_),
    .ZN(_05250_));
 NOR2_X1 _28293_ (.A1(net94),
    .A2(_05096_),
    .ZN(_05251_));
 AOI21_X1 _28294_ (.A(_04864_),
    .B1(_05017_),
    .B2(_04993_),
    .ZN(_05252_));
 OAI21_X1 _28295_ (.A(_04931_),
    .B1(_05251_),
    .B2(_05252_),
    .ZN(_05253_));
 NOR2_X1 _28296_ (.A1(_04987_),
    .A2(_05010_),
    .ZN(_05254_));
 OR3_X1 _28297_ (.A1(_04930_),
    .A2(_05030_),
    .A3(_05254_),
    .ZN(_05255_));
 AOI221_X2 _28298_ (.A(_04920_),
    .B1(_04997_),
    .B2(_05250_),
    .C1(_05253_),
    .C2(_05255_),
    .ZN(_05256_));
 NAND3_X1 _28299_ (.A1(_04899_),
    .A2(_05132_),
    .A3(_05106_),
    .ZN(_05257_));
 OAI21_X1 _28300_ (.A(_05224_),
    .B1(_05018_),
    .B2(_05008_),
    .ZN(_05258_));
 OAI21_X1 _28301_ (.A(_05257_),
    .B1(_05258_),
    .B2(_04983_),
    .ZN(_05259_));
 OAI21_X1 _28302_ (.A(_05078_),
    .B1(_05067_),
    .B2(_15274_),
    .ZN(_05260_));
 OAI21_X1 _28303_ (.A(_04966_),
    .B1(_05067_),
    .B2(net819),
    .ZN(_05261_));
 MUX2_X1 _28304_ (.A(_05260_),
    .B(_05261_),
    .S(_04970_),
    .Z(_05262_));
 MUX2_X1 _28305_ (.A(_05259_),
    .B(_05262_),
    .S(_04932_),
    .Z(_05263_));
 AOI211_X2 _28306_ (.A(_05037_),
    .B(_05256_),
    .C1(_05263_),
    .C2(_05075_),
    .ZN(_05264_));
 NOR2_X1 _28307_ (.A1(net1156),
    .A2(_05044_),
    .ZN(_05265_));
 OAI21_X1 _28308_ (.A(_04930_),
    .B1(_04881_),
    .B2(_04864_),
    .ZN(_05266_));
 AOI221_X2 _28309_ (.A(_04920_),
    .B1(_05265_),
    .B2(_05266_),
    .C1(_04975_),
    .C2(_04865_),
    .ZN(_05267_));
 NOR2_X1 _28310_ (.A1(_04991_),
    .A2(_05192_),
    .ZN(_05268_));
 NOR3_X4 _28311_ (.A1(_05092_),
    .A2(_04940_),
    .A3(_04946_),
    .ZN(_05269_));
 NOR2_X2 _28312_ (.A1(_05269_),
    .A2(_04956_),
    .ZN(_05270_));
 OAI221_X2 _28313_ (.A(_05268_),
    .B1(_05270_),
    .B2(_04983_),
    .C1(net97),
    .C2(_05083_),
    .ZN(_05271_));
 NOR2_X1 _28314_ (.A1(_05039_),
    .A2(_04960_),
    .ZN(_05272_));
 OAI21_X1 _28315_ (.A(_04992_),
    .B1(_05096_),
    .B2(_05272_),
    .ZN(_05273_));
 AND3_X2 _28316_ (.A1(_05267_),
    .A2(_05271_),
    .A3(_05273_),
    .ZN(_05274_));
 OAI22_X1 _28317_ (.A1(_05071_),
    .A2(_04947_),
    .B1(_05011_),
    .B2(net1155),
    .ZN(_05275_));
 OAI21_X4 _28318_ (.A(_04901_),
    .B1(_04958_),
    .B2(_04959_),
    .ZN(_05276_));
 OAI22_X1 _28319_ (.A1(_04998_),
    .A2(_04993_),
    .B1(_05276_),
    .B2(_05105_),
    .ZN(_05277_));
 AOI21_X1 _28320_ (.A(_05275_),
    .B1(_05277_),
    .B2(_15264_),
    .ZN(_05278_));
 NOR2_X1 _28321_ (.A1(_04933_),
    .A2(_05278_),
    .ZN(_05279_));
 AOI21_X1 _28322_ (.A(_05105_),
    .B1(_05049_),
    .B2(_05224_),
    .ZN(_05280_));
 NOR2_X1 _28323_ (.A1(net1153),
    .A2(_05276_),
    .ZN(_05281_));
 NOR4_X1 _28324_ (.A1(_04978_),
    .A2(_05265_),
    .A3(_05280_),
    .A4(_05281_),
    .ZN(_05282_));
 NOR4_X1 _28325_ (.A1(_05274_),
    .A2(_05006_),
    .A3(_05279_),
    .A4(_05282_),
    .ZN(_05283_));
 NAND2_X1 _28326_ (.A1(_15268_),
    .A2(_04970_),
    .ZN(_05284_));
 NAND4_X1 _28327_ (.A1(_05064_),
    .A2(_05068_),
    .A3(_05028_),
    .A4(_05284_),
    .ZN(_05285_));
 AOI21_X1 _28328_ (.A(_04991_),
    .B1(_04975_),
    .B2(net189),
    .ZN(_05286_));
 NAND2_X1 _28329_ (.A1(_05285_),
    .A2(_05286_),
    .ZN(_05287_));
 NAND3_X1 _28330_ (.A1(_04983_),
    .A2(_05064_),
    .A3(_04986_),
    .ZN(_05288_));
 NAND3_X1 _28331_ (.A1(_05105_),
    .A2(_04921_),
    .A3(_05068_),
    .ZN(_05289_));
 AOI21_X1 _28332_ (.A(_04973_),
    .B1(_05288_),
    .B2(_05289_),
    .ZN(_05290_));
 OAI22_X1 _28333_ (.A1(_05127_),
    .A2(_04993_),
    .B1(_05084_),
    .B2(_05023_),
    .ZN(_05291_));
 OAI221_X1 _28334_ (.A(_05088_),
    .B1(_05287_),
    .B2(_05290_),
    .C1(_05291_),
    .C2(_04933_),
    .ZN(_05292_));
 AOI21_X1 _28335_ (.A(_05019_),
    .B1(_05222_),
    .B2(_05051_),
    .ZN(_05293_));
 INV_X1 _28336_ (.A(_15274_),
    .ZN(_05294_));
 NAND2_X1 _28337_ (.A1(_05294_),
    .A2(_04898_),
    .ZN(_05295_));
 AOI21_X1 _28338_ (.A(_04982_),
    .B1(_05293_),
    .B2(_05295_),
    .ZN(_05296_));
 MUX2_X1 _28339_ (.A(net1155),
    .B(_15267_),
    .S(_04971_),
    .Z(_05297_));
 AOI21_X2 _28340_ (.A(_04980_),
    .B1(_05079_),
    .B2(_05297_),
    .ZN(_05298_));
 AOI21_X1 _28341_ (.A(_05292_),
    .B1(_05296_),
    .B2(_05298_),
    .ZN(_05299_));
 NAND2_X1 _28342_ (.A1(_05143_),
    .A2(_05005_),
    .ZN(_05300_));
 AOI21_X1 _28343_ (.A(_04901_),
    .B1(_04902_),
    .B2(_04965_),
    .ZN(_05301_));
 OR4_X1 _28344_ (.A1(_04977_),
    .A2(_05046_),
    .A3(_05254_),
    .A4(_05301_),
    .ZN(_05302_));
 AOI21_X4 _28345_ (.A(_04901_),
    .B1(_05041_),
    .B2(_05042_),
    .ZN(_05303_));
 OR2_X1 _28346_ (.A1(_04902_),
    .A2(_05177_),
    .ZN(_05304_));
 AOI21_X4 _28347_ (.A(_05023_),
    .B1(_04952_),
    .B2(_04955_),
    .ZN(_05305_));
 NOR2_X1 _28348_ (.A1(_05305_),
    .A2(_05269_),
    .ZN(_05306_));
 OAI221_X1 _28349_ (.A(_04981_),
    .B1(_05303_),
    .B2(_05304_),
    .C1(_05306_),
    .C2(_04899_),
    .ZN(_05307_));
 AOI21_X2 _28350_ (.A(_05064_),
    .B1(_05302_),
    .B2(_05307_),
    .ZN(_05308_));
 NOR2_X1 _28351_ (.A1(_05294_),
    .A2(_04904_),
    .ZN(_05309_));
 NOR2_X1 _28352_ (.A1(_15270_),
    .A2(_04896_),
    .ZN(_05310_));
 AOI221_X1 _28353_ (.A(_05310_),
    .B1(_04955_),
    .B2(_04952_),
    .C1(_04902_),
    .C2(_05222_),
    .ZN(_05311_));
 OAI33_X1 _28354_ (.A1(_05030_),
    .A2(_05160_),
    .A3(_05309_),
    .B1(_05311_),
    .B2(_05144_),
    .B3(_04981_),
    .ZN(_05312_));
 AOI211_X2 _28355_ (.A(_05300_),
    .B(_05308_),
    .C1(_05312_),
    .C2(_05101_),
    .ZN(_05313_));
 OR4_X2 _28356_ (.A1(_05283_),
    .A2(_05264_),
    .A3(_05299_),
    .A4(_05313_),
    .ZN(_00147_));
 OAI22_X1 _28357_ (.A1(_15267_),
    .A2(_05044_),
    .B1(_05177_),
    .B2(_05051_),
    .ZN(_05314_));
 AOI21_X1 _28358_ (.A(_05004_),
    .B1(_05111_),
    .B2(_05314_),
    .ZN(_05315_));
 NAND2_X1 _28359_ (.A1(_05008_),
    .A2(_15276_),
    .ZN(_05316_));
 OAI221_X1 _28360_ (.A(_05155_),
    .B1(_05316_),
    .B2(_05127_),
    .C1(_04947_),
    .C2(net1113),
    .ZN(_05317_));
 OAI21_X1 _28361_ (.A(_05315_),
    .B1(_05317_),
    .B2(_05114_),
    .ZN(_05318_));
 AND2_X1 _28362_ (.A1(_04935_),
    .A2(_04905_),
    .ZN(_05319_));
 OAI21_X1 _28363_ (.A(_05079_),
    .B1(_05319_),
    .B2(_05243_),
    .ZN(_05320_));
 NAND3_X1 _28364_ (.A1(_05087_),
    .A2(_04994_),
    .A3(_05320_),
    .ZN(_05321_));
 NOR2_X1 _28365_ (.A1(_05051_),
    .A2(_05056_),
    .ZN(_05322_));
 OAI21_X1 _28366_ (.A(_05322_),
    .B1(_05125_),
    .B2(_05014_),
    .ZN(_05323_));
 AND3_X1 _28367_ (.A1(_05075_),
    .A2(_05321_),
    .A3(_05323_),
    .ZN(_05324_));
 OAI21_X1 _28368_ (.A(_05005_),
    .B1(_05318_),
    .B2(_05324_),
    .ZN(_05325_));
 NAND2_X1 _28369_ (.A1(_04971_),
    .A2(_05116_),
    .ZN(_05326_));
 OAI221_X1 _28370_ (.A(_05056_),
    .B1(_05148_),
    .B2(_05326_),
    .C1(_05061_),
    .C2(_15258_),
    .ZN(_05327_));
 OAI21_X1 _28371_ (.A(_05059_),
    .B1(_05014_),
    .B2(_04983_),
    .ZN(_05328_));
 NOR2_X1 _28372_ (.A1(_04992_),
    .A2(_05328_),
    .ZN(_05329_));
 NOR2_X1 _28373_ (.A1(_05101_),
    .A2(_05329_),
    .ZN(_05330_));
 NAND2_X1 _28374_ (.A1(_04932_),
    .A2(_05191_),
    .ZN(_05331_));
 AOI21_X1 _28375_ (.A(_15264_),
    .B1(_05248_),
    .B2(_05331_),
    .ZN(_05332_));
 NAND2_X1 _28376_ (.A1(net159),
    .A2(_04931_),
    .ZN(_05333_));
 OAI221_X1 _28377_ (.A(_05127_),
    .B1(_05164_),
    .B2(_05009_),
    .C1(_05333_),
    .C2(_04900_),
    .ZN(_05334_));
 AOI21_X1 _28378_ (.A(net94),
    .B1(_15258_),
    .B2(_05217_),
    .ZN(_05335_));
 OR3_X1 _28379_ (.A1(_04998_),
    .A2(_05030_),
    .A3(_05335_),
    .ZN(_05336_));
 AOI21_X1 _28380_ (.A(_05332_),
    .B1(_05334_),
    .B2(_05336_),
    .ZN(_05337_));
 AOI221_X1 _28381_ (.A(_05143_),
    .B1(_05327_),
    .B2(_05330_),
    .C1(_05337_),
    .C2(_05065_),
    .ZN(_05338_));
 OAI21_X1 _28382_ (.A(_05170_),
    .B1(_04900_),
    .B2(net188),
    .ZN(_05339_));
 OAI21_X1 _28383_ (.A(_05004_),
    .B1(_05339_),
    .B2(_04978_),
    .ZN(_05340_));
 OAI21_X1 _28384_ (.A(_05047_),
    .B1(_04996_),
    .B2(_05019_),
    .ZN(_05341_));
 NOR2_X1 _28385_ (.A1(_04956_),
    .A2(_05177_),
    .ZN(_05342_));
 NAND2_X1 _28386_ (.A1(_04900_),
    .A2(_05342_),
    .ZN(_05343_));
 NAND2_X1 _28387_ (.A1(_04864_),
    .A2(_04901_),
    .ZN(_05344_));
 AOI221_X2 _28388_ (.A(_04931_),
    .B1(_04975_),
    .B2(_05344_),
    .C1(_05199_),
    .C2(net818),
    .ZN(_05345_));
 AOI21_X1 _28389_ (.A(_04980_),
    .B1(_05343_),
    .B2(_05345_),
    .ZN(_05346_));
 AOI21_X1 _28390_ (.A(_04933_),
    .B1(_05058_),
    .B2(_05127_),
    .ZN(_05347_));
 NOR3_X1 _28391_ (.A1(_05051_),
    .A2(_05305_),
    .A3(_05269_),
    .ZN(_05348_));
 AOI21_X1 _28392_ (.A(_05348_),
    .B1(_05177_),
    .B2(_15276_),
    .ZN(_05349_));
 AOI221_X2 _28393_ (.A(_05340_),
    .B1(_05341_),
    .B2(_05346_),
    .C1(_05347_),
    .C2(_05349_),
    .ZN(_05350_));
 INV_X1 _28394_ (.A(_15272_),
    .ZN(_05351_));
 MUX2_X1 _28395_ (.A(_05351_),
    .B(_05027_),
    .S(_04997_),
    .Z(_05352_));
 AOI22_X2 _28396_ (.A1(net95),
    .A2(_04975_),
    .B1(_05059_),
    .B2(_04971_),
    .ZN(_05353_));
 NOR3_X4 _28397_ (.A1(_04881_),
    .A2(_04940_),
    .A3(_04946_),
    .ZN(_05354_));
 AOI21_X1 _28398_ (.A(_04932_),
    .B1(_05354_),
    .B2(_15264_),
    .ZN(_05355_));
 AOI221_X2 _28399_ (.A(_05101_),
    .B1(_05352_),
    .B2(_04992_),
    .C1(_05353_),
    .C2(_05355_),
    .ZN(_05356_));
 AOI21_X1 _28400_ (.A(_05061_),
    .B1(_04966_),
    .B2(_05276_),
    .ZN(_05357_));
 OAI22_X1 _28401_ (.A1(net96),
    .A2(_05132_),
    .B1(_05083_),
    .B2(_05023_),
    .ZN(_05358_));
 AOI21_X1 _28402_ (.A(_04900_),
    .B1(_05048_),
    .B2(_05049_),
    .ZN(_05359_));
 OAI22_X1 _28403_ (.A1(_05008_),
    .A2(_05011_),
    .B1(_05276_),
    .B2(_15264_),
    .ZN(_05360_));
 NAND2_X1 _28404_ (.A1(_05064_),
    .A2(_04992_),
    .ZN(_05361_));
 OAI33_X1 _28405_ (.A1(_05114_),
    .A2(_05357_),
    .A3(_05358_),
    .B1(_05359_),
    .B2(_05360_),
    .B3(_05361_),
    .ZN(_05362_));
 OAI21_X1 _28406_ (.A(_05143_),
    .B1(_05356_),
    .B2(_05362_),
    .ZN(_05363_));
 NAND2_X1 _28407_ (.A1(_04915_),
    .A2(_05363_),
    .ZN(_05364_));
 OAI22_X1 _28408_ (.A1(_05325_),
    .A2(_05338_),
    .B1(_05350_),
    .B2(_05364_),
    .ZN(_00148_));
 NAND3_X1 _28409_ (.A1(_05051_),
    .A2(_04966_),
    .A3(_05106_),
    .ZN(_05365_));
 OAI221_X1 _28410_ (.A(_04971_),
    .B1(_04998_),
    .B2(net898),
    .C1(_05276_),
    .C2(net1153),
    .ZN(_05366_));
 NAND3_X1 _28411_ (.A1(_04982_),
    .A2(_05365_),
    .A3(_05366_),
    .ZN(_05367_));
 OAI22_X1 _28412_ (.A1(_15267_),
    .A2(_05154_),
    .B1(_04993_),
    .B2(_04998_),
    .ZN(_05368_));
 NAND2_X1 _28413_ (.A1(_05056_),
    .A2(_05368_),
    .ZN(_05369_));
 AOI21_X1 _28414_ (.A(_05004_),
    .B1(_05367_),
    .B2(_05369_),
    .ZN(_05370_));
 OAI21_X1 _28415_ (.A(_05018_),
    .B1(_05058_),
    .B2(_05310_),
    .ZN(_05371_));
 NAND2_X1 _28416_ (.A1(net896),
    .A2(_04903_),
    .ZN(_05372_));
 AOI21_X1 _28417_ (.A(_04931_),
    .B1(_05013_),
    .B2(_05372_),
    .ZN(_05373_));
 NAND3_X1 _28418_ (.A1(_04970_),
    .A2(_04966_),
    .A3(_04968_),
    .ZN(_05374_));
 AND2_X1 _28419_ (.A1(_05015_),
    .A2(_05374_),
    .ZN(_05375_));
 AOI221_X2 _28420_ (.A(_05143_),
    .B1(_05371_),
    .B2(_05373_),
    .C1(_05375_),
    .C2(_04932_),
    .ZN(_05376_));
 NOR4_X1 _28421_ (.A1(_05065_),
    .A2(_04915_),
    .A3(_05370_),
    .A4(_05376_),
    .ZN(_05377_));
 NAND2_X1 _28422_ (.A1(_05064_),
    .A2(_04909_),
    .ZN(_05378_));
 OAI21_X1 _28423_ (.A(_05043_),
    .B1(_05281_),
    .B2(_04904_),
    .ZN(_05379_));
 NAND2_X1 _28424_ (.A1(_05038_),
    .A2(_05379_),
    .ZN(_05380_));
 AOI22_X1 _28425_ (.A1(_04881_),
    .A2(_05228_),
    .B1(_05306_),
    .B2(_04903_),
    .ZN(_05381_));
 AOI21_X1 _28426_ (.A(_04915_),
    .B1(_05381_),
    .B2(_04991_),
    .ZN(_05382_));
 AOI21_X1 _28427_ (.A(_04903_),
    .B1(_05048_),
    .B2(_05115_),
    .ZN(_05383_));
 AOI21_X1 _28428_ (.A(_05383_),
    .B1(_05199_),
    .B2(net94),
    .ZN(_05384_));
 NOR2_X1 _28429_ (.A1(_04973_),
    .A2(_04947_),
    .ZN(_05385_));
 OAI21_X1 _28430_ (.A(_05200_),
    .B1(_05067_),
    .B2(_05007_),
    .ZN(_05386_));
 AOI21_X1 _28431_ (.A(_05385_),
    .B1(_05386_),
    .B2(_04899_),
    .ZN(_05387_));
 MUX2_X1 _28432_ (.A(_05384_),
    .B(_05387_),
    .S(_04991_),
    .Z(_05388_));
 AOI221_X2 _28433_ (.A(_05378_),
    .B1(_05382_),
    .B2(_05380_),
    .C1(_05388_),
    .C2(_04915_),
    .ZN(_05389_));
 AND3_X2 _28434_ (.A1(_04902_),
    .A2(_05078_),
    .A3(_05106_),
    .ZN(_05390_));
 AOI21_X1 _28435_ (.A(_05177_),
    .B1(_04985_),
    .B2(_15268_),
    .ZN(_05391_));
 AOI21_X2 _28436_ (.A(_05390_),
    .B1(_05391_),
    .B2(_04970_),
    .ZN(_05392_));
 OR2_X2 _28437_ (.A1(_05392_),
    .A2(_04991_),
    .ZN(_05393_));
 NAND3_X1 _28438_ (.A1(net159),
    .A2(_05017_),
    .A3(_05030_),
    .ZN(_05394_));
 NAND3_X1 _28439_ (.A1(_04931_),
    .A2(_05231_),
    .A3(_05394_),
    .ZN(_05395_));
 AND2_X1 _28440_ (.A1(_05064_),
    .A2(_05395_),
    .ZN(_05396_));
 AOI221_X1 _28441_ (.A(_04977_),
    .B1(_05154_),
    .B2(_05147_),
    .C1(_05222_),
    .C2(_04974_),
    .ZN(_05397_));
 MUX2_X1 _28442_ (.A(_05020_),
    .B(_05295_),
    .S(_04997_),
    .Z(_05398_));
 AOI21_X1 _28443_ (.A(_05397_),
    .B1(_05398_),
    .B2(_05038_),
    .ZN(_05399_));
 AOI221_X1 _28444_ (.A(_05198_),
    .B1(_05393_),
    .B2(_05396_),
    .C1(_05399_),
    .C2(_04980_),
    .ZN(_05400_));
 NOR2_X1 _28445_ (.A1(_05143_),
    .A2(_05005_),
    .ZN(_05401_));
 OAI22_X1 _28446_ (.A1(_15267_),
    .A2(_05044_),
    .B1(_05083_),
    .B2(_05071_),
    .ZN(_05402_));
 NAND2_X1 _28447_ (.A1(_04982_),
    .A2(_05402_),
    .ZN(_05403_));
 NAND3_X1 _28448_ (.A1(_05075_),
    .A2(_05401_),
    .A3(_05403_),
    .ZN(_05404_));
 AND3_X1 _28449_ (.A1(_05038_),
    .A2(_05154_),
    .A3(_04915_),
    .ZN(_05405_));
 AOI21_X1 _28450_ (.A(_04986_),
    .B1(_04914_),
    .B2(_04991_),
    .ZN(_05406_));
 AOI21_X1 _28451_ (.A(_04899_),
    .B1(_04991_),
    .B2(_04914_),
    .ZN(_05407_));
 OAI22_X1 _28452_ (.A1(_15264_),
    .A2(_05406_),
    .B1(_05407_),
    .B2(_05068_),
    .ZN(_05408_));
 NAND3_X1 _28453_ (.A1(_04981_),
    .A2(_04915_),
    .A3(_05284_),
    .ZN(_05409_));
 AOI21_X1 _28454_ (.A(_05199_),
    .B1(_05409_),
    .B2(_04998_),
    .ZN(_05410_));
 OAI33_X1 _28455_ (.A1(_15258_),
    .A2(_05405_),
    .A3(_05408_),
    .B1(_05410_),
    .B2(_04859_),
    .B3(_04862_),
    .ZN(_05411_));
 OAI21_X1 _28456_ (.A(_05019_),
    .B1(_05030_),
    .B2(_05020_),
    .ZN(_05412_));
 NAND3_X1 _28457_ (.A1(_04992_),
    .A2(_04994_),
    .A3(_05412_),
    .ZN(_05413_));
 MUX2_X1 _28458_ (.A(_05076_),
    .B(_05391_),
    .S(_04971_),
    .Z(_05414_));
 OAI21_X1 _28459_ (.A(_05413_),
    .B1(_05056_),
    .B2(_05414_),
    .ZN(_05415_));
 NAND2_X1 _28460_ (.A1(_05065_),
    .A2(_04916_),
    .ZN(_05416_));
 OAI22_X1 _28461_ (.A1(_05404_),
    .A2(_05411_),
    .B1(_05415_),
    .B2(_05416_),
    .ZN(_05417_));
 OR4_X2 _28462_ (.A1(_05417_),
    .A2(_05389_),
    .A3(_05400_),
    .A4(_05377_),
    .ZN(_00149_));
 OAI221_X2 _28463_ (.A(_05143_),
    .B1(_05203_),
    .B2(_05075_),
    .C1(_04925_),
    .C2(net1152),
    .ZN(_05418_));
 AOI21_X1 _28464_ (.A(_05065_),
    .B1(_05127_),
    .B2(_15278_),
    .ZN(_05419_));
 NAND2_X1 _28465_ (.A1(net188),
    .A2(_15283_),
    .ZN(_05420_));
 NAND3_X1 _28466_ (.A1(_05079_),
    .A2(_05028_),
    .A3(_05420_),
    .ZN(_05421_));
 AOI21_X1 _28467_ (.A(_05418_),
    .B1(_05419_),
    .B2(_05421_),
    .ZN(_05422_));
 MUX2_X1 _28468_ (.A(_05023_),
    .B(net160),
    .S(_05018_),
    .Z(_05423_));
 AOI22_X2 _28469_ (.A1(net96),
    .A2(_04975_),
    .B1(_05423_),
    .B2(_04900_),
    .ZN(_05424_));
 NOR3_X1 _28470_ (.A1(_05004_),
    .A2(_05114_),
    .A3(_05424_),
    .ZN(_05425_));
 AOI21_X1 _28471_ (.A(_04905_),
    .B1(_04968_),
    .B2(_05132_),
    .ZN(_05426_));
 NOR4_X1 _28472_ (.A1(_04978_),
    .A2(_05004_),
    .A3(_05385_),
    .A4(_05426_),
    .ZN(_05427_));
 OR3_X1 _28473_ (.A1(_05005_),
    .A2(_05425_),
    .A3(_05427_),
    .ZN(_05428_));
 NOR2_X1 _28474_ (.A1(_05105_),
    .A2(_05344_),
    .ZN(_05429_));
 OAI21_X1 _28475_ (.A(_05018_),
    .B1(_04899_),
    .B2(_04973_),
    .ZN(_05430_));
 OAI221_X2 _28476_ (.A(_04921_),
    .B1(_05429_),
    .B2(_05430_),
    .C1(_05019_),
    .C2(_15279_),
    .ZN(_05431_));
 AOI21_X1 _28477_ (.A(_05067_),
    .B1(_04993_),
    .B2(net159),
    .ZN(_05432_));
 NOR3_X1 _28478_ (.A1(_04921_),
    .A2(_05082_),
    .A3(_05432_),
    .ZN(_05433_));
 NOR2_X1 _28479_ (.A1(_04992_),
    .A2(_05433_),
    .ZN(_05434_));
 NOR3_X1 _28480_ (.A1(_04983_),
    .A2(_04956_),
    .A3(_05269_),
    .ZN(_05435_));
 AOI221_X1 _28481_ (.A(_04902_),
    .B1(_05017_),
    .B2(_05000_),
    .C1(_05191_),
    .C2(net159),
    .ZN(_05436_));
 NOR3_X1 _28482_ (.A1(_05101_),
    .A2(_05435_),
    .A3(_05436_),
    .ZN(_05437_));
 AOI221_X1 _28483_ (.A(_04898_),
    .B1(_05017_),
    .B2(_05222_),
    .C1(_05191_),
    .C2(_04864_),
    .ZN(_05438_));
 NOR3_X1 _28484_ (.A1(_04904_),
    .A2(_05303_),
    .A3(_05269_),
    .ZN(_05439_));
 NOR3_X1 _28485_ (.A1(_04921_),
    .A2(_05438_),
    .A3(_05439_),
    .ZN(_05440_));
 NOR2_X1 _28486_ (.A1(_05437_),
    .A2(_05440_),
    .ZN(_05441_));
 AOI221_X2 _28487_ (.A(_05143_),
    .B1(_05431_),
    .B2(_05434_),
    .C1(_05441_),
    .C2(_05056_),
    .ZN(_05442_));
 OAI21_X1 _28488_ (.A(_05059_),
    .B1(_04997_),
    .B2(_05008_),
    .ZN(_05443_));
 NAND2_X1 _28489_ (.A1(_04904_),
    .A2(_05443_),
    .ZN(_05444_));
 AOI21_X1 _28490_ (.A(_05063_),
    .B1(_05228_),
    .B2(net189),
    .ZN(_05445_));
 NOR2_X1 _28491_ (.A1(_05305_),
    .A2(_05354_),
    .ZN(_05446_));
 MUX2_X1 _28492_ (.A(net1156),
    .B(_05222_),
    .S(_04985_),
    .Z(_05447_));
 MUX2_X1 _28493_ (.A(_05446_),
    .B(_05447_),
    .S(_04970_),
    .Z(_05448_));
 AOI221_X2 _28494_ (.A(_04932_),
    .B1(_05444_),
    .B2(_05445_),
    .C1(_05448_),
    .C2(_05064_),
    .ZN(_05449_));
 OAI21_X1 _28495_ (.A(_04986_),
    .B1(_15258_),
    .B2(_04987_),
    .ZN(_05450_));
 AND3_X1 _28496_ (.A1(_04900_),
    .A2(_05450_),
    .A3(_05183_),
    .ZN(_05451_));
 NAND2_X1 _28497_ (.A1(_04905_),
    .A2(_05200_),
    .ZN(_05452_));
 NOR2_X1 _28498_ (.A1(_05069_),
    .A2(_05452_),
    .ZN(_05453_));
 NOR3_X1 _28499_ (.A1(_05361_),
    .A2(_05451_),
    .A3(_05453_),
    .ZN(_05454_));
 AOI21_X2 _28500_ (.A(_05450_),
    .B1(_05051_),
    .B2(net96),
    .ZN(_05455_));
 NOR3_X1 _28501_ (.A1(_15277_),
    .A2(_15286_),
    .A3(_04998_),
    .ZN(_05456_));
 NOR3_X1 _28502_ (.A1(_04933_),
    .A2(_05455_),
    .A3(_05456_),
    .ZN(_05457_));
 NOR4_X1 _28503_ (.A1(_05143_),
    .A2(_05449_),
    .A3(_05454_),
    .A4(_05457_),
    .ZN(_05458_));
 NAND3_X1 _28504_ (.A1(_04904_),
    .A2(_04931_),
    .A3(_04997_),
    .ZN(_05459_));
 NAND3_X1 _28505_ (.A1(_15267_),
    .A2(_05164_),
    .A3(_05459_),
    .ZN(_05460_));
 NAND2_X1 _28506_ (.A1(_05294_),
    .A2(net94),
    .ZN(_05461_));
 OAI21_X1 _28507_ (.A(_05333_),
    .B1(_05461_),
    .B2(_05248_),
    .ZN(_05462_));
 OAI21_X1 _28508_ (.A(_05460_),
    .B1(_05462_),
    .B2(_15267_),
    .ZN(_05463_));
 NOR2_X1 _28509_ (.A1(_04864_),
    .A2(_04930_),
    .ZN(_05464_));
 OAI21_X1 _28510_ (.A(_05028_),
    .B1(_04930_),
    .B2(_04901_),
    .ZN(_05465_));
 OR2_X1 _28511_ (.A1(_04930_),
    .A2(net708),
    .ZN(_05466_));
 AOI221_X2 _28512_ (.A(_05063_),
    .B1(_05191_),
    .B2(_05464_),
    .C1(_05465_),
    .C2(_05466_),
    .ZN(_05467_));
 NAND3_X1 _28513_ (.A1(_04931_),
    .A2(_05059_),
    .A3(_05078_),
    .ZN(_05468_));
 NAND3_X1 _28514_ (.A1(_05105_),
    .A2(_05160_),
    .A3(_05468_),
    .ZN(_05469_));
 AOI21_X1 _28515_ (.A(_05464_),
    .B1(_05191_),
    .B2(_04991_),
    .ZN(_05470_));
 OAI221_X2 _28516_ (.A(_05469_),
    .B1(_05470_),
    .B2(_04905_),
    .C1(_15258_),
    .C2(_05160_),
    .ZN(_05471_));
 AOI221_X2 _28517_ (.A(_05004_),
    .B1(_05463_),
    .B2(_05467_),
    .C1(_05471_),
    .C2(_05065_),
    .ZN(_05472_));
 OAI33_X1 _28518_ (.A1(_05422_),
    .A2(_05428_),
    .A3(_05442_),
    .B1(_05458_),
    .B2(_05472_),
    .B3(_04915_),
    .ZN(_00150_));
 AOI21_X1 _28519_ (.A(_05056_),
    .B1(_04975_),
    .B2(_05008_),
    .ZN(_05473_));
 AOI21_X1 _28520_ (.A(_05354_),
    .B1(_05303_),
    .B2(_05061_),
    .ZN(_05474_));
 OAI221_X1 _28521_ (.A(_05473_),
    .B1(_05474_),
    .B2(net96),
    .C1(_15267_),
    .C2(_05011_),
    .ZN(_05475_));
 OAI221_X1 _28522_ (.A(_05087_),
    .B1(_05083_),
    .B2(net188),
    .C1(_05342_),
    .C2(_15283_),
    .ZN(_05476_));
 NAND3_X1 _28523_ (.A1(_05075_),
    .A2(_05475_),
    .A3(_05476_),
    .ZN(_05477_));
 NAND3_X1 _28524_ (.A1(_15276_),
    .A2(_05049_),
    .A3(_05200_),
    .ZN(_05478_));
 OAI21_X1 _28525_ (.A(_05478_),
    .B1(_05184_),
    .B2(_15276_),
    .ZN(_05479_));
 OAI21_X1 _28526_ (.A(_05027_),
    .B1(_05061_),
    .B2(_05294_),
    .ZN(_05480_));
 AOI21_X1 _28527_ (.A(_05087_),
    .B1(_05127_),
    .B2(_05480_),
    .ZN(_05481_));
 AOI22_X1 _28528_ (.A1(_05111_),
    .A2(_05479_),
    .B1(_05481_),
    .B2(_05298_),
    .ZN(_05482_));
 NAND3_X1 _28529_ (.A1(_04916_),
    .A2(_05477_),
    .A3(_05482_),
    .ZN(_05483_));
 OAI21_X1 _28530_ (.A(_04966_),
    .B1(_04947_),
    .B2(_05222_),
    .ZN(_05484_));
 OR2_X1 _28531_ (.A1(_05305_),
    .A2(_05354_),
    .ZN(_05485_));
 AOI21_X2 _28532_ (.A(_05484_),
    .B1(_05485_),
    .B2(_15283_),
    .ZN(_05486_));
 AOI21_X1 _28533_ (.A(_15276_),
    .B1(_05102_),
    .B2(_05231_),
    .ZN(_05487_));
 OR2_X1 _28534_ (.A1(_04982_),
    .A2(_05117_),
    .ZN(_05488_));
 OAI221_X2 _28535_ (.A(_05075_),
    .B1(_05087_),
    .B2(_05486_),
    .C1(_05487_),
    .C2(_05488_),
    .ZN(_05489_));
 NOR2_X1 _28536_ (.A1(_05008_),
    .A2(_05061_),
    .ZN(_05490_));
 AOI21_X1 _28537_ (.A(_05014_),
    .B1(_05127_),
    .B2(_15264_),
    .ZN(_05491_));
 AOI21_X1 _28538_ (.A(_05490_),
    .B1(_05491_),
    .B2(_15283_),
    .ZN(_05492_));
 OAI21_X1 _28539_ (.A(_04982_),
    .B1(_05127_),
    .B2(net1113),
    .ZN(_05493_));
 OAI221_X2 _28540_ (.A(_05065_),
    .B1(_04982_),
    .B2(_05492_),
    .C1(_05493_),
    .C2(_05455_),
    .ZN(_05494_));
 NAND4_X2 _28541_ (.A1(_05004_),
    .A2(_05005_),
    .A3(_05489_),
    .A4(_05494_),
    .ZN(_05495_));
 NOR3_X1 _28542_ (.A1(_04932_),
    .A2(_05068_),
    .A3(_05057_),
    .ZN(_05496_));
 OAI21_X1 _28543_ (.A(_05011_),
    .B1(_05019_),
    .B2(_05038_),
    .ZN(_05497_));
 AOI21_X1 _28544_ (.A(_05496_),
    .B1(_05497_),
    .B2(_15267_),
    .ZN(_05498_));
 OAI221_X1 _28545_ (.A(_05217_),
    .B1(_05498_),
    .B2(net96),
    .C1(_05044_),
    .C2(net1157),
    .ZN(_05499_));
 OR3_X1 _28546_ (.A1(_05075_),
    .A2(_05198_),
    .A3(_05499_),
    .ZN(_05500_));
 AND2_X1 _28547_ (.A1(_15264_),
    .A2(_05354_),
    .ZN(_05501_));
 AOI21_X1 _28548_ (.A(_15264_),
    .B1(_05011_),
    .B2(_05049_),
    .ZN(_05502_));
 OAI21_X2 _28549_ (.A(_05087_),
    .B1(_05501_),
    .B2(_05502_),
    .ZN(_05503_));
 AOI21_X1 _28550_ (.A(_04960_),
    .B1(_04975_),
    .B2(_15258_),
    .ZN(_05504_));
 AOI21_X2 _28551_ (.A(_05228_),
    .B1(_05030_),
    .B2(_05079_),
    .ZN(_05505_));
 OAI221_X2 _28552_ (.A(_05503_),
    .B1(_05504_),
    .B2(_05087_),
    .C1(net96),
    .C2(_05505_),
    .ZN(_05506_));
 NOR2_X1 _28553_ (.A1(_05065_),
    .A2(_05198_),
    .ZN(_05507_));
 AOI22_X4 _28554_ (.A1(_05105_),
    .A2(_04935_),
    .B1(_05041_),
    .B2(_05042_),
    .ZN(_05508_));
 AOI22_X4 _28555_ (.A1(_05154_),
    .A2(_04993_),
    .B1(_05508_),
    .B2(_04996_),
    .ZN(_05509_));
 NAND4_X1 _28556_ (.A1(net189),
    .A2(_04971_),
    .A3(_05041_),
    .A4(_05042_),
    .ZN(_05510_));
 OAI21_X1 _28557_ (.A(_05510_),
    .B1(_05019_),
    .B2(_15272_),
    .ZN(_05511_));
 AOI22_X4 _28558_ (.A1(_05509_),
    .A2(_05176_),
    .B1(_05511_),
    .B2(_05187_),
    .ZN(_05512_));
 NOR3_X1 _28559_ (.A1(_05243_),
    .A2(_05024_),
    .A3(_04998_),
    .ZN(_05513_));
 NOR2_X1 _28560_ (.A1(_15286_),
    .A2(_05019_),
    .ZN(_05514_));
 OR2_X1 _28561_ (.A1(_05513_),
    .A2(_05514_),
    .ZN(_05515_));
 OAI21_X4 _28562_ (.A(_05106_),
    .B1(_05127_),
    .B2(net96),
    .ZN(_05516_));
 AOI21_X2 _28563_ (.A(_05133_),
    .B1(_15276_),
    .B2(_05516_),
    .ZN(_05517_));
 OAI221_X2 _28564_ (.A(_05512_),
    .B1(_05515_),
    .B2(_05361_),
    .C1(_05114_),
    .C2(_05517_),
    .ZN(_05518_));
 AOI22_X2 _28565_ (.A1(_05506_),
    .A2(_05507_),
    .B1(_05518_),
    .B2(_05401_),
    .ZN(_05519_));
 NAND4_X4 _28566_ (.A1(_05519_),
    .A2(_05495_),
    .A3(_05500_),
    .A4(_05483_),
    .ZN(_00151_));
 INV_X1 _28567_ (.A(net1017),
    .ZN(_05520_));
 NOR2_X1 _28568_ (.A1(_05520_),
    .A2(_09102_),
    .ZN(_05521_));
 NOR2_X1 _28569_ (.A1(net1017),
    .A2(_11841_),
    .ZN(_05522_));
 XNOR2_X2 _28570_ (.A(_11184_),
    .B(_11119_),
    .ZN(_05523_));
 XNOR2_X2 _28571_ (.A(_11122_),
    .B(_05523_),
    .ZN(_05524_));
 XNOR2_X2 _28572_ (.A(_13842_),
    .B(_11166_),
    .ZN(_05525_));
 XNOR2_X2 _28573_ (.A(_05525_),
    .B(_05524_),
    .ZN(_05526_));
 MUX2_X2 _28574_ (.A(_05521_),
    .B(_05522_),
    .S(_05526_),
    .Z(_05527_));
 OR3_X2 _28575_ (.A1(net1017),
    .A2(_09074_),
    .A3(_00405_),
    .ZN(_05528_));
 NAND3_X2 _28576_ (.A1(net1017),
    .A2(_11938_),
    .A3(_00405_),
    .ZN(_05529_));
 NAND2_X4 _28577_ (.A1(_05528_),
    .A2(_05529_),
    .ZN(_05530_));
 NOR2_X4 _28578_ (.A1(_05530_),
    .A2(_05527_),
    .ZN(_05531_));
 INV_X4 _28579_ (.A(_05531_),
    .ZN(_05532_));
 BUF_X16 _28580_ (.A(_05532_),
    .Z(_05533_));
 BUF_X32 _28581_ (.A(_05533_),
    .Z(_05534_));
 BUF_X32 _28582_ (.A(_05534_),
    .Z(_15296_));
 XNOR2_X1 _28583_ (.A(\sa03_sr[0] ),
    .B(net661),
    .ZN(_05535_));
 NAND3_X1 _28584_ (.A1(net1019),
    .A2(_09856_),
    .A3(_11144_),
    .ZN(_05536_));
 NOR2_X1 _28585_ (.A1(net1019),
    .A2(_08973_),
    .ZN(_05537_));
 NAND2_X1 _28586_ (.A1(net966),
    .A2(_05537_),
    .ZN(_05538_));
 AOI21_X1 _28587_ (.A(_05535_),
    .B1(_05536_),
    .B2(_05538_),
    .ZN(_05539_));
 XOR2_X1 _28588_ (.A(\sa03_sr[0] ),
    .B(net661),
    .Z(_05540_));
 NAND2_X1 _28589_ (.A1(_11144_),
    .A2(_05537_),
    .ZN(_05541_));
 NAND3_X1 _28590_ (.A1(net1021),
    .A2(_09100_),
    .A3(net966),
    .ZN(_05542_));
 AOI21_X1 _28591_ (.A(_05540_),
    .B1(_05541_),
    .B2(_05542_),
    .ZN(_05543_));
 INV_X1 _28592_ (.A(net1019),
    .ZN(_05544_));
 NAND3_X1 _28593_ (.A1(_05544_),
    .A2(_09102_),
    .A3(_00406_),
    .ZN(_05545_));
 NAND2_X1 _28594_ (.A1(net1019),
    .A2(_11841_),
    .ZN(_05546_));
 OAI21_X1 _28595_ (.A(_05545_),
    .B1(_05546_),
    .B2(_00406_),
    .ZN(_05547_));
 OR3_X4 _28596_ (.A1(_05543_),
    .A2(_05539_),
    .A3(_05547_),
    .ZN(_05548_));
 INV_X8 _28597_ (.A(_05548_),
    .ZN(_05549_));
 BUF_X1 rebuffer495 (.A(_13835_),
    .Z(net958));
 BUF_X8 _28599_ (.A(_05549_),
    .Z(_15299_));
 XNOR2_X1 _28600_ (.A(_11219_),
    .B(_02927_),
    .ZN(_05551_));
 NAND3_X1 _28601_ (.A1(_06354_),
    .A2(net947),
    .A3(_11162_),
    .ZN(_05552_));
 NOR2_X1 _28602_ (.A1(_06354_),
    .A2(_08992_),
    .ZN(_05553_));
 NAND2_X1 _28603_ (.A1(_11160_),
    .A2(_05553_),
    .ZN(_05554_));
 AOI21_X2 _28604_ (.A(_05551_),
    .B1(_05552_),
    .B2(_05554_),
    .ZN(_05555_));
 XOR2_X1 _28605_ (.A(_11219_),
    .B(_02927_),
    .Z(_05556_));
 NAND2_X1 _28606_ (.A1(_11162_),
    .A2(_05553_),
    .ZN(_05557_));
 NAND3_X1 _28607_ (.A1(_06354_),
    .A2(_09022_),
    .A3(_11160_),
    .ZN(_05558_));
 AOI21_X2 _28608_ (.A(_05556_),
    .B1(_05557_),
    .B2(_05558_),
    .ZN(_05559_));
 NAND3_X1 _28609_ (.A1(_06367_),
    .A2(_09726_),
    .A3(_00407_),
    .ZN(_05560_));
 NAND2_X1 _28610_ (.A1(_06354_),
    .A2(_09726_),
    .ZN(_05561_));
 OAI21_X2 _28611_ (.A(_05560_),
    .B1(_05561_),
    .B2(_00407_),
    .ZN(_05562_));
 NOR3_X4 _28612_ (.A1(_05555_),
    .A2(_05559_),
    .A3(_05562_),
    .ZN(_05563_));
 INV_X8 _28613_ (.A(_05563_),
    .ZN(_05564_));
 BUF_X4 _28614_ (.A(_05564_),
    .Z(_05565_));
 BUF_X4 _28615_ (.A(_05565_),
    .Z(_05566_));
 BUF_X4 _28616_ (.A(_05566_),
    .Z(_15315_));
 BUF_X16 _28617_ (.A(_05548_),
    .Z(_05567_));
 BUF_X8 _28618_ (.A(_05567_),
    .Z(_15290_));
 BUF_X4 _28619_ (.A(_05563_),
    .Z(_05568_));
 BUF_X4 _28620_ (.A(_05568_),
    .Z(_05569_));
 BUF_X4 _28621_ (.A(_05569_),
    .Z(_05570_));
 BUF_X4 _28622_ (.A(_05570_),
    .Z(_15308_));
 XNOR2_X1 _28623_ (.A(_11202_),
    .B(_11187_),
    .ZN(_05571_));
 XNOR2_X1 _28624_ (.A(_11200_),
    .B(_05571_),
    .ZN(_05572_));
 XNOR2_X1 _28625_ (.A(_11262_),
    .B(_05572_),
    .ZN(_05573_));
 MUX2_X2 _28626_ (.A(\text_in_r[6] ),
    .B(_05573_),
    .S(net951),
    .Z(_05574_));
 XNOR2_X1 _28627_ (.A(_06430_),
    .B(_05574_),
    .ZN(_05575_));
 BUF_X4 _28628_ (.A(_05575_),
    .Z(_05576_));
 XNOR2_X1 _28629_ (.A(_11121_),
    .B(_13904_),
    .ZN(_05577_));
 XNOR2_X1 _28630_ (.A(_11183_),
    .B(_05577_),
    .ZN(_05578_));
 MUX2_X2 _28631_ (.A(\text_in_r[7] ),
    .B(_05578_),
    .S(_11207_),
    .Z(_05579_));
 XOR2_X2 _28632_ (.A(\u0.tmp_w[7] ),
    .B(_05579_),
    .Z(_05580_));
 BUF_X4 _28633_ (.A(_05580_),
    .Z(_05581_));
 OR2_X2 _28634_ (.A1(_05576_),
    .A2(_05581_),
    .ZN(_05582_));
 OR2_X1 _28635_ (.A1(_11191_),
    .A2(\text_in_r[4] ),
    .ZN(_05583_));
 XNOR2_X2 _28636_ (.A(_11248_),
    .B(_03011_),
    .ZN(_05584_));
 OAI211_X4 _28637_ (.A(_06407_),
    .B(_05583_),
    .C1(_05584_),
    .C2(_09824_),
    .ZN(_05585_));
 INV_X1 _28638_ (.A(_06407_),
    .ZN(_05586_));
 NAND2_X1 _28639_ (.A1(_09180_),
    .A2(\text_in_r[4] ),
    .ZN(_05587_));
 XOR2_X2 _28640_ (.A(_11248_),
    .B(_03011_),
    .Z(_05588_));
 OAI211_X4 _28641_ (.A(_05586_),
    .B(_05587_),
    .C1(_05588_),
    .C2(_09824_),
    .ZN(_05589_));
 AND2_X1 _28642_ (.A1(_05585_),
    .A2(_05589_),
    .ZN(_05590_));
 BUF_X4 _28643_ (.A(_05590_),
    .Z(_05591_));
 NOR2_X4 _28644_ (.A1(_05548_),
    .A2(_05564_),
    .ZN(_05592_));
 NAND2_X1 _28645_ (.A1(_05533_),
    .A2(_05592_),
    .ZN(_05593_));
 INV_X1 _28646_ (.A(\text_in_r[3] ),
    .ZN(_05594_));
 NAND2_X1 _28647_ (.A1(net582),
    .A2(_05594_),
    .ZN(_05595_));
 XNOR2_X2 _28648_ (.A(_11222_),
    .B(_02987_),
    .ZN(_05596_));
 OAI211_X4 _28649_ (.A(_06393_),
    .B(_05595_),
    .C1(_05596_),
    .C2(_08996_),
    .ZN(_05597_));
 BUF_X8 _28650_ (.A(_05597_),
    .Z(_05598_));
 INV_X1 _28651_ (.A(_06393_),
    .ZN(_05599_));
 NAND2_X1 _28652_ (.A1(net582),
    .A2(\text_in_r[3] ),
    .ZN(_05600_));
 XOR2_X2 _28653_ (.A(_11222_),
    .B(_02987_),
    .Z(_05601_));
 OAI211_X4 _28654_ (.A(_05599_),
    .B(_05600_),
    .C1(_05601_),
    .C2(_09135_),
    .ZN(_05602_));
 BUF_X8 _28655_ (.A(_05602_),
    .Z(_05603_));
 NAND2_X4 _28656_ (.A1(_05598_),
    .A2(_05603_),
    .ZN(_05604_));
 NOR2_X1 _28657_ (.A1(_05549_),
    .A2(_05568_),
    .ZN(_05605_));
 NOR2_X2 _28658_ (.A1(_05604_),
    .A2(_05605_),
    .ZN(_05606_));
 AOI21_X4 _28659_ (.A(_05591_),
    .B1(_05593_),
    .B2(_05606_),
    .ZN(_05607_));
 INV_X1 _28660_ (.A(_06416_),
    .ZN(_05608_));
 XNOR2_X1 _28661_ (.A(_11265_),
    .B(_11261_),
    .ZN(_05609_));
 NOR3_X1 _28662_ (.A1(_05608_),
    .A2(_08975_),
    .A3(_05609_),
    .ZN(_05610_));
 NOR3_X1 _28663_ (.A1(_06416_),
    .A2(_08975_),
    .A3(_05609_),
    .ZN(_05611_));
 MUX2_X2 _28664_ (.A(_05610_),
    .B(_05611_),
    .S(_03020_),
    .Z(_05612_));
 XOR2_X1 _28665_ (.A(_11265_),
    .B(_11261_),
    .Z(_05613_));
 NOR3_X1 _28666_ (.A1(_06416_),
    .A2(_00991_),
    .A3(_05613_),
    .ZN(_05614_));
 NOR3_X1 _28667_ (.A1(_05608_),
    .A2(_00991_),
    .A3(_05613_),
    .ZN(_05615_));
 MUX2_X1 _28668_ (.A(_05614_),
    .B(_05615_),
    .S(_03020_),
    .Z(_05616_));
 NAND3_X1 _28669_ (.A1(_06416_),
    .A2(_09135_),
    .A3(\text_in_r[5] ),
    .ZN(_05617_));
 NAND2_X1 _28670_ (.A1(_05608_),
    .A2(_09135_),
    .ZN(_05618_));
 OAI21_X2 _28671_ (.A(_05617_),
    .B1(_05618_),
    .B2(\text_in_r[5] ),
    .ZN(_05619_));
 NOR3_X4 _28672_ (.A1(_05612_),
    .A2(_05616_),
    .A3(_05619_),
    .ZN(_05620_));
 BUF_X4 _28673_ (.A(_05620_),
    .Z(_05621_));
 BUF_X4 _28674_ (.A(_05621_),
    .Z(_05622_));
 BUF_X4 _28675_ (.A(_05564_),
    .Z(_05623_));
 BUF_X4 _28676_ (.A(_05623_),
    .Z(_05624_));
 OAI21_X2 _28677_ (.A(_05624_),
    .B1(_05530_),
    .B2(_05527_),
    .ZN(_05625_));
 NOR2_X1 _28678_ (.A1(_09194_),
    .A2(\text_in_r[3] ),
    .ZN(_05626_));
 AOI211_X4 _28679_ (.A(_05599_),
    .B(_05626_),
    .C1(_05601_),
    .C2(_09075_),
    .ZN(_05627_));
 NOR2_X1 _28680_ (.A1(_09194_),
    .A2(_05594_),
    .ZN(_05628_));
 AOI211_X4 _28681_ (.A(_06393_),
    .B(_05628_),
    .C1(_05596_),
    .C2(net1085),
    .ZN(_05629_));
 NOR2_X2 _28682_ (.A1(_05627_),
    .A2(_05629_),
    .ZN(_05630_));
 BUF_X4 _28683_ (.A(_05630_),
    .Z(_05631_));
 BUF_X4 _28684_ (.A(_05631_),
    .Z(_05632_));
 CLKBUF_X3 _28685_ (.A(_05568_),
    .Z(_05633_));
 BUF_X4 _28686_ (.A(_15294_),
    .Z(_05634_));
 INV_X1 _28687_ (.A(_05634_),
    .ZN(_05635_));
 AOI21_X1 _28688_ (.A(_05632_),
    .B1(_05633_),
    .B2(_05635_),
    .ZN(_05636_));
 AOI21_X1 _28689_ (.A(_05622_),
    .B1(_05625_),
    .B2(_05636_),
    .ZN(_05637_));
 OR3_X2 _28690_ (.A1(_05612_),
    .A2(_05616_),
    .A3(_05619_),
    .ZN(_05638_));
 BUF_X4 _28691_ (.A(_05638_),
    .Z(_05639_));
 NOR2_X2 _28692_ (.A1(_05639_),
    .A2(_05591_),
    .ZN(_05640_));
 INV_X2 clone106 (.A(net111),
    .ZN(net106));
 BUF_X4 _28694_ (.A(_15297_),
    .Z(_05642_));
 NAND3_X2 _28695_ (.A1(_05563_),
    .A2(_05598_),
    .A3(_05603_),
    .ZN(_05643_));
 BUF_X4 _28696_ (.A(_05643_),
    .Z(_05644_));
 NAND2_X1 _28697_ (.A1(_05567_),
    .A2(_05623_),
    .ZN(_05645_));
 NOR2_X1 _28698_ (.A1(_05532_),
    .A2(_05604_),
    .ZN(_05646_));
 OAI22_X1 _28699_ (.A1(net654),
    .A2(_05644_),
    .B1(_05645_),
    .B2(_05646_),
    .ZN(_05647_));
 AOI221_X1 _28700_ (.A(_05582_),
    .B1(_05607_),
    .B2(_05637_),
    .C1(_05640_),
    .C2(_05647_),
    .ZN(_05648_));
 BUF_X4 _28701_ (.A(_05639_),
    .Z(_05649_));
 CLKBUF_X3 _28702_ (.A(_05649_),
    .Z(_05650_));
 NOR2_X1 _28703_ (.A1(_05534_),
    .A2(_05632_),
    .ZN(_05651_));
 BUF_X8 clone14 (.A(_07377_),
    .Z(net14));
 BUF_X4 _28705_ (.A(_05598_),
    .Z(_05653_));
 BUF_X8 _28706_ (.A(_05603_),
    .Z(_05654_));
 NAND3_X2 _28707_ (.A1(_15306_),
    .A2(_05653_),
    .A3(_05654_),
    .ZN(_05655_));
 BUF_X4 _28708_ (.A(_05627_),
    .Z(_05656_));
 BUF_X8 _28709_ (.A(_05629_),
    .Z(_05657_));
 OAI22_X4 _28710_ (.A1(net526),
    .A2(_05530_),
    .B1(_05656_),
    .B2(_05657_),
    .ZN(_05658_));
 NAND2_X1 _28711_ (.A1(_05655_),
    .A2(_05658_),
    .ZN(_05659_));
 OAI221_X1 _28712_ (.A(_05650_),
    .B1(_05651_),
    .B2(_05645_),
    .C1(_05659_),
    .C2(_15315_),
    .ZN(_05660_));
 AOI21_X4 _28713_ (.A(_05567_),
    .B1(_05598_),
    .B2(_05603_),
    .ZN(_05661_));
 NOR3_X4 _28714_ (.A1(_05564_),
    .A2(_05627_),
    .A3(_05629_),
    .ZN(_05662_));
 BUF_X4 _28715_ (.A(_15293_),
    .Z(_05663_));
 BUF_X8 _28716_ (.A(_05663_),
    .Z(_05664_));
 BUF_X4 _28717_ (.A(_05633_),
    .Z(_05665_));
 NOR3_X4 _28718_ (.A1(net909),
    .A2(_05627_),
    .A3(_05629_),
    .ZN(_05666_));
 NOR2_X1 _28719_ (.A1(_05665_),
    .A2(_05666_),
    .ZN(_05667_));
 AOI221_X1 _28720_ (.A(_05661_),
    .B1(_05662_),
    .B2(net902),
    .C1(_05658_),
    .C2(_05667_),
    .ZN(_05668_));
 OAI21_X1 _28721_ (.A(_05660_),
    .B1(_05668_),
    .B2(_05650_),
    .ZN(_05669_));
 NAND2_X4 _28722_ (.A1(_05585_),
    .A2(_05589_),
    .ZN(_05670_));
 BUF_X4 _28723_ (.A(_05670_),
    .Z(_05671_));
 BUF_X4 _28724_ (.A(_05671_),
    .Z(_05672_));
 BUF_X4 _28725_ (.A(_05672_),
    .Z(_05673_));
 OAI21_X1 _28726_ (.A(_05648_),
    .B1(_05669_),
    .B2(_05673_),
    .ZN(_05674_));
 XOR2_X2 _28727_ (.A(_06430_),
    .B(_05574_),
    .Z(_05675_));
 BUF_X4 _28728_ (.A(_05675_),
    .Z(_05676_));
 OR2_X2 _28729_ (.A1(_05676_),
    .A2(_05581_),
    .ZN(_05677_));
 BUF_X8 clone108 (.A(net934),
    .Z(net108));
 NOR3_X4 _28731_ (.A1(_05563_),
    .A2(_05627_),
    .A3(_05629_),
    .ZN(_05679_));
 OAI21_X4 _28732_ (.A(_05563_),
    .B1(_05627_),
    .B2(_05629_),
    .ZN(_05680_));
 AOI21_X2 _28733_ (.A(_05680_),
    .B1(_05622_),
    .B2(_05664_),
    .ZN(_05681_));
 OAI21_X2 _28734_ (.A(_15292_),
    .B1(_05681_),
    .B2(_05679_),
    .ZN(_05682_));
 BUF_X4 _28735_ (.A(_15300_),
    .Z(_05683_));
 INV_X2 _28736_ (.A(_05683_),
    .ZN(_05684_));
 NOR2_X1 _28737_ (.A1(_05684_),
    .A2(_05621_),
    .ZN(_05685_));
 AND2_X1 _28738_ (.A1(_05528_),
    .A2(_05529_),
    .ZN(_05686_));
 NAND2_X1 _28739_ (.A1(net1017),
    .A2(_10571_),
    .ZN(_05687_));
 NAND2_X1 _28740_ (.A1(_05520_),
    .A2(_10571_),
    .ZN(_05688_));
 MUX2_X2 _28741_ (.A(_05687_),
    .B(_05688_),
    .S(_05526_),
    .Z(_05689_));
 AOI21_X4 _28742_ (.A(_05548_),
    .B1(_05686_),
    .B2(_05689_),
    .ZN(_05690_));
 AOI21_X1 _28743_ (.A(_05685_),
    .B1(_05690_),
    .B2(_05622_),
    .ZN(_05691_));
 OAI21_X4 _28744_ (.A(_05623_),
    .B1(_05656_),
    .B2(_05657_),
    .ZN(_05692_));
 BUF_X4 _28745_ (.A(_05639_),
    .Z(_05693_));
 NAND3_X2 _28746_ (.A1(_05683_),
    .A2(_05653_),
    .A3(_05654_),
    .ZN(_05694_));
 NOR2_X1 _28747_ (.A1(_05693_),
    .A2(_05694_),
    .ZN(_05695_));
 BUF_X4 _28748_ (.A(_05631_),
    .Z(_05696_));
 XNOR2_X1 _28749_ (.A(_05639_),
    .B(_05696_),
    .ZN(_05697_));
 INV_X8 _28750_ (.A(_05663_),
    .ZN(_05698_));
 AOI21_X1 _28751_ (.A(_05695_),
    .B1(_05697_),
    .B2(_05698_),
    .ZN(_05699_));
 OAI221_X1 _28752_ (.A(_05682_),
    .B1(_05691_),
    .B2(_05692_),
    .C1(_15315_),
    .C2(_05699_),
    .ZN(_05700_));
 CLKBUF_X3 _28753_ (.A(_05696_),
    .Z(_05701_));
 NAND2_X1 _28754_ (.A1(_05565_),
    .A2(_05639_),
    .ZN(_05702_));
 CLKBUF_X3 _28755_ (.A(_05592_),
    .Z(_05703_));
 BUF_X4 _28756_ (.A(_05531_),
    .Z(_05704_));
 AOI21_X1 _28757_ (.A(_05703_),
    .B1(_15290_),
    .B2(_05704_),
    .ZN(_05705_));
 OAI221_X1 _28758_ (.A(_05701_),
    .B1(_05702_),
    .B2(net902),
    .C1(_05705_),
    .C2(_05693_),
    .ZN(_05706_));
 NAND3_X1 _28759_ (.A1(_05664_),
    .A2(_05570_),
    .A3(_05693_),
    .ZN(_05707_));
 AOI21_X1 _28760_ (.A(_05624_),
    .B1(_05622_),
    .B2(_15290_),
    .ZN(_05708_));
 BUF_X8 _28761_ (.A(_05531_),
    .Z(_05709_));
 BUF_X16 _28762_ (.A(_05709_),
    .Z(_15291_));
 NAND2_X1 _28763_ (.A1(_15299_),
    .A2(_05566_),
    .ZN(_05710_));
 OAI221_X1 _28764_ (.A(_05707_),
    .B1(_05708_),
    .B2(net105),
    .C1(_05649_),
    .C2(_05710_),
    .ZN(_05711_));
 OAI21_X1 _28765_ (.A(_05706_),
    .B1(_05711_),
    .B2(_05701_),
    .ZN(_05712_));
 BUF_X4 _28766_ (.A(_05591_),
    .Z(_05713_));
 BUF_X4 _28767_ (.A(_05713_),
    .Z(_05714_));
 BUF_X4 _28768_ (.A(_05714_),
    .Z(_05715_));
 MUX2_X1 _28769_ (.A(_05700_),
    .B(_05712_),
    .S(_05715_),
    .Z(_05716_));
 BUF_X4 _28770_ (.A(_05591_),
    .Z(_05717_));
 CLKBUF_X3 _28771_ (.A(_05717_),
    .Z(_05718_));
 BUF_X4 _28772_ (.A(_05604_),
    .Z(_05719_));
 BUF_X4 _28773_ (.A(_05719_),
    .Z(_05720_));
 OAI21_X2 _28774_ (.A(net910),
    .B1(_05656_),
    .B2(_05657_),
    .ZN(_05721_));
 OAI221_X2 _28775_ (.A(_05665_),
    .B1(_05720_),
    .B2(_05634_),
    .C1(_05721_),
    .C2(_05704_),
    .ZN(_05722_));
 AOI21_X2 _28776_ (.A(_05563_),
    .B1(_05653_),
    .B2(_05654_),
    .ZN(_05723_));
 BUF_X4 _28777_ (.A(_05723_),
    .Z(_05724_));
 NAND2_X1 _28778_ (.A1(_05684_),
    .A2(_05724_),
    .ZN(_05725_));
 AND3_X1 _28779_ (.A1(_05718_),
    .A2(_05722_),
    .A3(_05725_),
    .ZN(_05726_));
 BUF_X4 _28780_ (.A(_15302_),
    .Z(_05727_));
 BUF_X4 _28781_ (.A(_05727_),
    .Z(_05728_));
 OAI21_X4 _28782_ (.A(_05548_),
    .B1(_05530_),
    .B2(net527),
    .ZN(_05729_));
 MUX2_X1 _28783_ (.A(_05634_),
    .B(_05729_),
    .S(_05631_),
    .Z(_05730_));
 AOI221_X1 _28784_ (.A(_05717_),
    .B1(_05679_),
    .B2(_05728_),
    .C1(_05730_),
    .C2(_05665_),
    .ZN(_05731_));
 NOR3_X1 _28785_ (.A1(_05650_),
    .A2(_05726_),
    .A3(_05731_),
    .ZN(_05732_));
 CLKBUF_X3 _28786_ (.A(_05621_),
    .Z(_05733_));
 BUF_X4 _28787_ (.A(_05604_),
    .Z(_05734_));
 MUX2_X1 _28788_ (.A(_15297_),
    .B(_05729_),
    .S(_05568_),
    .Z(_05735_));
 AOI21_X4 _28789_ (.A(_05713_),
    .B1(_05734_),
    .B2(_05735_),
    .ZN(_05736_));
 NOR2_X1 _28790_ (.A1(_15292_),
    .A2(_05643_),
    .ZN(_05737_));
 NAND3_X4 _28791_ (.A1(_05549_),
    .A2(_05598_),
    .A3(_05603_),
    .ZN(_05738_));
 OAI21_X1 _28792_ (.A(_05738_),
    .B1(_05632_),
    .B2(_05635_),
    .ZN(_05739_));
 BUF_X4 _28793_ (.A(_05565_),
    .Z(_05740_));
 AOI21_X1 _28794_ (.A(_05737_),
    .B1(_05739_),
    .B2(_05740_),
    .ZN(_05741_));
 BUF_X4 _28795_ (.A(_05632_),
    .Z(_05742_));
 AOI22_X1 _28796_ (.A1(_15313_),
    .A2(_05742_),
    .B1(_05724_),
    .B2(net902),
    .ZN(_05743_));
 AOI221_X1 _28797_ (.A(_05733_),
    .B1(_05736_),
    .B2(_05741_),
    .C1(_05743_),
    .C2(_05718_),
    .ZN(_05744_));
 NOR3_X2 _28798_ (.A1(_05744_),
    .A2(_05732_),
    .A3(_05676_),
    .ZN(_05745_));
 BUF_X4 _28799_ (.A(_05581_),
    .Z(_05746_));
 NOR2_X1 _28800_ (.A1(_05576_),
    .A2(_05649_),
    .ZN(_05747_));
 BUF_X4 _28801_ (.A(_05719_),
    .Z(_05748_));
 NAND2_X1 _28802_ (.A1(_05634_),
    .A2(_05748_),
    .ZN(_05749_));
 NAND3_X4 _28803_ (.A1(_15297_),
    .A2(_05653_),
    .A3(_05654_),
    .ZN(_05750_));
 AND3_X1 _28804_ (.A1(_15308_),
    .A2(_05749_),
    .A3(_05750_),
    .ZN(_05751_));
 INV_X1 _28805_ (.A(_15292_),
    .ZN(_05752_));
 OAI21_X1 _28806_ (.A(_05718_),
    .B1(_05692_),
    .B2(_05752_),
    .ZN(_05753_));
 NOR3_X4 _28807_ (.A1(_05567_),
    .A2(_05627_),
    .A3(_05629_),
    .ZN(_05754_));
 BUF_X4 _28808_ (.A(_05734_),
    .Z(_05755_));
 AOI21_X1 _28809_ (.A(_05754_),
    .B1(_05755_),
    .B2(_15291_),
    .ZN(_05756_));
 AOI21_X4 _28810_ (.A(_05663_),
    .B1(_05653_),
    .B2(_05654_),
    .ZN(_05757_));
 AOI21_X1 _28811_ (.A(_05757_),
    .B1(_05742_),
    .B2(_05684_),
    .ZN(_05758_));
 CLKBUF_X3 _28812_ (.A(_05624_),
    .Z(_05759_));
 MUX2_X1 _28813_ (.A(_05756_),
    .B(_05758_),
    .S(_05759_),
    .Z(_05760_));
 OAI221_X1 _28814_ (.A(_05747_),
    .B1(_05751_),
    .B2(_05753_),
    .C1(_05760_),
    .C2(_05715_),
    .ZN(_05761_));
 NOR2_X1 _28815_ (.A1(_05576_),
    .A2(_05733_),
    .ZN(_05762_));
 NAND2_X1 _28816_ (.A1(net910),
    .A2(_05670_),
    .ZN(_05763_));
 NOR2_X1 _28817_ (.A1(_05755_),
    .A2(_05763_),
    .ZN(_05764_));
 AOI21_X4 _28818_ (.A(net655),
    .B1(_05653_),
    .B2(_05654_),
    .ZN(_05765_));
 OR2_X1 _28819_ (.A1(_15308_),
    .A2(_05765_),
    .ZN(_05766_));
 NAND3_X2 _28820_ (.A1(net102),
    .A2(_05653_),
    .A3(_05654_),
    .ZN(_05767_));
 OAI21_X1 _28821_ (.A(_05728_),
    .B1(_05656_),
    .B2(_05657_),
    .ZN(_05768_));
 AOI21_X1 _28822_ (.A(_05759_),
    .B1(_05767_),
    .B2(_05768_),
    .ZN(_05769_));
 NOR2_X1 _28823_ (.A1(_05673_),
    .A2(_05769_),
    .ZN(_05770_));
 OAI221_X1 _28824_ (.A(_05762_),
    .B1(_05764_),
    .B2(_05766_),
    .C1(_05770_),
    .C2(_05607_),
    .ZN(_05771_));
 NAND3_X1 _28825_ (.A1(_05746_),
    .A2(_05761_),
    .A3(_05771_),
    .ZN(_05772_));
 OAI221_X2 _28826_ (.A(_05674_),
    .B1(_05716_),
    .B2(_05677_),
    .C1(_05745_),
    .C2(_05772_),
    .ZN(_00152_));
 OAI21_X4 _28827_ (.A(net1028),
    .B1(_05627_),
    .B2(_05629_),
    .ZN(_05773_));
 NOR3_X4 _28828_ (.A1(_05627_),
    .A2(_05663_),
    .A3(_05629_),
    .ZN(_05774_));
 NOR2_X2 _28829_ (.A1(_05565_),
    .A2(_05774_),
    .ZN(_05775_));
 OAI22_X4 _28830_ (.A1(_05634_),
    .A2(_05632_),
    .B1(_05738_),
    .B2(net508),
    .ZN(_05776_));
 AOI221_X2 _28831_ (.A(_05671_),
    .B1(_05775_),
    .B2(_05773_),
    .C1(_05776_),
    .C2(_05740_),
    .ZN(_05777_));
 OAI21_X2 _28832_ (.A(_05549_),
    .B1(_05656_),
    .B2(_05657_),
    .ZN(_05778_));
 OAI22_X1 _28833_ (.A1(net102),
    .A2(_05719_),
    .B1(_05778_),
    .B2(net100),
    .ZN(_05779_));
 AOI221_X1 _28834_ (.A(_05713_),
    .B1(_05724_),
    .B2(_15290_),
    .C1(_05779_),
    .C2(_05570_),
    .ZN(_05780_));
 NOR3_X1 _28835_ (.A1(_05733_),
    .A2(_05777_),
    .A3(_05780_),
    .ZN(_05781_));
 NAND2_X4 _28836_ (.A1(_05620_),
    .A2(_05671_),
    .ZN(_05782_));
 OAI21_X4 _28837_ (.A(_15292_),
    .B1(_05656_),
    .B2(_05657_),
    .ZN(_05783_));
 OAI21_X1 _28838_ (.A(_05783_),
    .B1(_05748_),
    .B2(_05534_),
    .ZN(_05784_));
 NOR2_X1 _28839_ (.A1(_15308_),
    .A2(_05784_),
    .ZN(_05785_));
 AOI21_X1 _28840_ (.A(_05759_),
    .B1(_05721_),
    .B2(_05750_),
    .ZN(_05786_));
 NAND2_X2 _28841_ (.A1(_05621_),
    .A2(_05713_),
    .ZN(_05787_));
 AOI21_X1 _28842_ (.A(_05665_),
    .B1(_05778_),
    .B2(_05767_),
    .ZN(_05788_));
 NOR3_X2 _28843_ (.A1(_05752_),
    .A2(_05656_),
    .A3(_05657_),
    .ZN(_05789_));
 OAI21_X2 _28844_ (.A(_05633_),
    .B1(_05632_),
    .B2(_05634_),
    .ZN(_05790_));
 NOR2_X1 _28845_ (.A1(_05789_),
    .A2(_05790_),
    .ZN(_05791_));
 OAI33_X1 _28846_ (.A1(_05782_),
    .A2(_05785_),
    .A3(_05786_),
    .B1(_05787_),
    .B2(_05788_),
    .B3(_05791_),
    .ZN(_05792_));
 OR3_X2 _28847_ (.A1(_05781_),
    .A2(_05746_),
    .A3(_05792_),
    .ZN(_05793_));
 OR2_X1 _28848_ (.A1(_05719_),
    .A2(_05690_),
    .ZN(_05794_));
 AOI21_X1 _28849_ (.A(_05774_),
    .B1(_05719_),
    .B2(_05642_),
    .ZN(_05795_));
 MUX2_X1 _28850_ (.A(_05794_),
    .B(_05795_),
    .S(_05633_),
    .Z(_05796_));
 NAND2_X1 _28851_ (.A1(_05581_),
    .A2(_05640_),
    .ZN(_05797_));
 OAI21_X1 _28852_ (.A(_05676_),
    .B1(_05796_),
    .B2(_05797_),
    .ZN(_05798_));
 AND2_X1 _28853_ (.A1(_05580_),
    .A2(_05621_),
    .ZN(_05799_));
 NAND2_X1 _28854_ (.A1(_05714_),
    .A2(_05799_),
    .ZN(_05800_));
 AOI21_X1 _28855_ (.A(_05800_),
    .B1(_05662_),
    .B2(net105),
    .ZN(_05801_));
 CLKBUF_X3 _28856_ (.A(_05633_),
    .Z(_05802_));
 NAND2_X1 _28857_ (.A1(_05534_),
    .A2(_05661_),
    .ZN(_05803_));
 NAND2_X1 _28858_ (.A1(_05802_),
    .A2(_05803_),
    .ZN(_05804_));
 NAND2_X1 _28859_ (.A1(_05655_),
    .A2(_05804_),
    .ZN(_05805_));
 NAND3_X1 _28860_ (.A1(_05633_),
    .A2(_05767_),
    .A3(_05783_),
    .ZN(_05806_));
 AND2_X1 _28861_ (.A1(_05778_),
    .A2(_05750_),
    .ZN(_05807_));
 OAI21_X1 _28862_ (.A(_05806_),
    .B1(_05807_),
    .B2(_05570_),
    .ZN(_05808_));
 OAI22_X1 _28863_ (.A1(_05698_),
    .A2(_05692_),
    .B1(_05738_),
    .B2(_05533_),
    .ZN(_05809_));
 NAND3_X4 _28864_ (.A1(_05564_),
    .A2(_05653_),
    .A3(_05654_),
    .ZN(_05810_));
 NAND2_X1 _28865_ (.A1(_05810_),
    .A2(_05680_),
    .ZN(_05811_));
 AOI21_X1 _28866_ (.A(_05809_),
    .B1(_05811_),
    .B2(_15290_),
    .ZN(_05812_));
 MUX2_X1 _28867_ (.A(_05808_),
    .B(_05812_),
    .S(_05672_),
    .Z(_05813_));
 NAND2_X2 _28868_ (.A1(_05580_),
    .A2(_05639_),
    .ZN(_05814_));
 INV_X1 _28869_ (.A(_05814_),
    .ZN(_05815_));
 AOI221_X2 _28870_ (.A(_05798_),
    .B1(_05801_),
    .B2(_05805_),
    .C1(_05813_),
    .C2(_05815_),
    .ZN(_05816_));
 NOR2_X2 _28871_ (.A1(_05698_),
    .A2(_05569_),
    .ZN(_05817_));
 INV_X1 _28872_ (.A(_15306_),
    .ZN(_05818_));
 NOR2_X1 _28873_ (.A1(_05818_),
    .A2(_05624_),
    .ZN(_05819_));
 OAI21_X1 _28874_ (.A(_05742_),
    .B1(_05817_),
    .B2(_05819_),
    .ZN(_05820_));
 AOI21_X4 _28875_ (.A(_05564_),
    .B1(_05598_),
    .B2(_05603_),
    .ZN(_05821_));
 NOR2_X2 _28876_ (.A1(_05679_),
    .A2(_05821_),
    .ZN(_05822_));
 OAI22_X1 _28877_ (.A1(net654),
    .A2(_05692_),
    .B1(_05822_),
    .B2(_05704_),
    .ZN(_05823_));
 AOI221_X2 _28878_ (.A(_05814_),
    .B1(_05820_),
    .B2(_05736_),
    .C1(_05823_),
    .C2(_05718_),
    .ZN(_05824_));
 NOR2_X2 _28879_ (.A1(_05765_),
    .A2(_05774_),
    .ZN(_05825_));
 OAI221_X1 _28880_ (.A(_05715_),
    .B1(_05692_),
    .B2(_15290_),
    .C1(_05825_),
    .C2(_15315_),
    .ZN(_05826_));
 OAI21_X1 _28881_ (.A(_05826_),
    .B1(_05662_),
    .B2(_05715_),
    .ZN(_05827_));
 NAND2_X1 _28882_ (.A1(_05580_),
    .A2(_05621_),
    .ZN(_05828_));
 OAI22_X1 _28883_ (.A1(_05566_),
    .A2(_05717_),
    .B1(_05810_),
    .B2(_05549_),
    .ZN(_05829_));
 NAND2_X1 _28884_ (.A1(_05704_),
    .A2(_05720_),
    .ZN(_05830_));
 NAND2_X1 _28885_ (.A1(_05740_),
    .A2(_05717_),
    .ZN(_05831_));
 OAI22_X2 _28886_ (.A1(_05714_),
    .A2(_05830_),
    .B1(_05831_),
    .B2(_05748_),
    .ZN(_05832_));
 AOI221_X2 _28887_ (.A(_05828_),
    .B1(_05829_),
    .B2(_15296_),
    .C1(_05832_),
    .C2(_15290_),
    .ZN(_05833_));
 AOI21_X1 _28888_ (.A(_05824_),
    .B1(_05827_),
    .B2(_05833_),
    .ZN(_05834_));
 OAI21_X1 _28889_ (.A(_05721_),
    .B1(_05738_),
    .B2(net103),
    .ZN(_05835_));
 AOI221_X1 _28890_ (.A(_05639_),
    .B1(_05724_),
    .B2(_15292_),
    .C1(_05835_),
    .C2(_05570_),
    .ZN(_05836_));
 AOI221_X1 _28891_ (.A(_05621_),
    .B1(_05703_),
    .B2(_05750_),
    .C1(_05724_),
    .C2(_05534_),
    .ZN(_05837_));
 OR3_X1 _28892_ (.A1(_05673_),
    .A2(_05836_),
    .A3(_05837_),
    .ZN(_05838_));
 NOR2_X1 _28893_ (.A1(net100),
    .A2(_05568_),
    .ZN(_05839_));
 NAND2_X1 _28894_ (.A1(_05693_),
    .A2(_05717_),
    .ZN(_05840_));
 INV_X1 _28895_ (.A(_05642_),
    .ZN(_05841_));
 NOR2_X1 _28896_ (.A1(_05841_),
    .A2(_05565_),
    .ZN(_05842_));
 NOR4_X2 _28897_ (.A1(_05842_),
    .A2(_05839_),
    .A3(_05840_),
    .A4(_05755_),
    .ZN(_05843_));
 OAI21_X1 _28898_ (.A(_05622_),
    .B1(_05742_),
    .B2(_15292_),
    .ZN(_05844_));
 NOR3_X1 _28899_ (.A1(_05729_),
    .A2(_05831_),
    .A3(_05844_),
    .ZN(_05845_));
 AOI221_X2 _28900_ (.A(_05630_),
    .B1(_05592_),
    .B2(_05532_),
    .C1(_05564_),
    .C2(_05683_),
    .ZN(_05846_));
 NOR3_X1 _28901_ (.A1(_15316_),
    .A2(_05622_),
    .A3(_05720_),
    .ZN(_05847_));
 NOR3_X1 _28902_ (.A1(_05718_),
    .A2(_05846_),
    .A3(_05847_),
    .ZN(_05848_));
 NOR4_X2 _28903_ (.A1(_05746_),
    .A2(_05843_),
    .A3(_05845_),
    .A4(_05848_),
    .ZN(_05849_));
 AOI21_X2 _28904_ (.A(_05676_),
    .B1(_05838_),
    .B2(_05849_),
    .ZN(_05850_));
 AOI22_X4 _28905_ (.A1(_05793_),
    .A2(_05816_),
    .B1(_05834_),
    .B2(_05850_),
    .ZN(_00153_));
 NAND2_X1 _28906_ (.A1(_05676_),
    .A2(_05581_),
    .ZN(_05851_));
 OAI211_X2 _28907_ (.A(_05802_),
    .B(_05694_),
    .C1(_05701_),
    .C2(_15296_),
    .ZN(_05852_));
 OAI21_X1 _28908_ (.A(_05783_),
    .B1(_05720_),
    .B2(_05664_),
    .ZN(_05853_));
 OAI211_X2 _28909_ (.A(_05649_),
    .B(_05852_),
    .C1(_05853_),
    .C2(_15308_),
    .ZN(_05854_));
 NOR3_X1 _28910_ (.A1(_05534_),
    .A2(_05719_),
    .A3(_05703_),
    .ZN(_05855_));
 OAI21_X1 _28911_ (.A(_05658_),
    .B1(_05569_),
    .B2(_05534_),
    .ZN(_05856_));
 NOR2_X2 _28912_ (.A1(net100),
    .A2(_05623_),
    .ZN(_05857_));
 AOI221_X2 _28913_ (.A(_05855_),
    .B1(_05856_),
    .B2(net902),
    .C1(_05738_),
    .C2(_05857_),
    .ZN(_05858_));
 OAI211_X2 _28914_ (.A(_05715_),
    .B(_05854_),
    .C1(_05858_),
    .C2(_05650_),
    .ZN(_05859_));
 NOR2_X1 _28915_ (.A1(_15296_),
    .A2(_15299_),
    .ZN(_05860_));
 NOR3_X1 _28916_ (.A1(_05755_),
    .A2(_05860_),
    .A3(_05857_),
    .ZN(_05861_));
 OAI21_X1 _28917_ (.A(_05649_),
    .B1(_05701_),
    .B2(_15316_),
    .ZN(_05862_));
 MUX2_X1 _28918_ (.A(net102),
    .B(_05729_),
    .S(_05569_),
    .Z(_05863_));
 MUX2_X1 _28919_ (.A(_15313_),
    .B(_05863_),
    .S(_05701_),
    .Z(_05864_));
 OAI221_X1 _28920_ (.A(_05673_),
    .B1(_05861_),
    .B2(_05862_),
    .C1(_05864_),
    .C2(_05650_),
    .ZN(_05865_));
 AND2_X1 _28921_ (.A1(_05859_),
    .A2(_05865_),
    .ZN(_05866_));
 AOI21_X4 _28922_ (.A(_05698_),
    .B1(_05597_),
    .B2(_05602_),
    .ZN(_05867_));
 OAI21_X4 _28923_ (.A(_05569_),
    .B1(_05867_),
    .B2(_05754_),
    .ZN(_05868_));
 NAND3_X1 _28924_ (.A1(_05635_),
    .A2(_05653_),
    .A3(_05654_),
    .ZN(_05869_));
 NAND3_X1 _28925_ (.A1(_05566_),
    .A2(_05658_),
    .A3(_05869_),
    .ZN(_05870_));
 AOI21_X2 _28926_ (.A(_05672_),
    .B1(_05868_),
    .B2(_05870_),
    .ZN(_05871_));
 NOR3_X4 _28927_ (.A1(_05549_),
    .A2(_05627_),
    .A3(_05629_),
    .ZN(_05872_));
 NOR2_X1 _28928_ (.A1(_05661_),
    .A2(_05872_),
    .ZN(_05873_));
 AOI221_X1 _28929_ (.A(_05713_),
    .B1(_05839_),
    .B2(_05873_),
    .C1(_05662_),
    .C2(_05818_),
    .ZN(_05874_));
 NOR4_X1 _28930_ (.A1(_05746_),
    .A2(_05649_),
    .A3(_05871_),
    .A4(_05874_),
    .ZN(_05875_));
 NOR2_X4 _28931_ (.A1(net659),
    .A2(_15294_),
    .ZN(_05876_));
 INV_X1 _28932_ (.A(_05876_),
    .ZN(_05877_));
 NOR2_X2 _28933_ (.A1(_05877_),
    .A2(_05643_),
    .ZN(_05878_));
 AOI221_X2 _28934_ (.A(_05878_),
    .B1(_05811_),
    .B2(_05690_),
    .C1(_05683_),
    .C2(_05724_),
    .ZN(_05879_));
 OAI221_X1 _28935_ (.A(_05799_),
    .B1(_05853_),
    .B2(_05759_),
    .C1(_05810_),
    .C2(_05841_),
    .ZN(_05880_));
 OAI221_X1 _28936_ (.A(_05576_),
    .B1(_05879_),
    .B2(_05800_),
    .C1(_05880_),
    .C2(_05715_),
    .ZN(_05881_));
 OR2_X2 _28937_ (.A1(_05875_),
    .A2(_05881_),
    .ZN(_05882_));
 BUF_X4 _28938_ (.A(_05671_),
    .Z(_05883_));
 OAI21_X1 _28939_ (.A(_05883_),
    .B1(_05748_),
    .B2(_05735_),
    .ZN(_05884_));
 NOR3_X1 _28940_ (.A1(_05742_),
    .A2(_05817_),
    .A3(_05857_),
    .ZN(_05885_));
 OR3_X1 _28941_ (.A1(_05746_),
    .A2(_05884_),
    .A3(_05885_),
    .ZN(_05886_));
 AOI22_X2 _28942_ (.A1(_05689_),
    .A2(_05686_),
    .B1(_05549_),
    .B2(_05565_),
    .ZN(_05887_));
 MUX2_X1 _28943_ (.A(_15311_),
    .B(_05887_),
    .S(_05713_),
    .Z(_05888_));
 NOR2_X1 _28944_ (.A1(_05755_),
    .A2(_05888_),
    .ZN(_05889_));
 NOR2_X1 _28945_ (.A1(_15320_),
    .A2(_05883_),
    .ZN(_05890_));
 NOR3_X1 _28946_ (.A1(_05570_),
    .A2(_05717_),
    .A3(_05729_),
    .ZN(_05891_));
 NOR3_X1 _28947_ (.A1(_05701_),
    .A2(_05890_),
    .A3(_05891_),
    .ZN(_05892_));
 OAI21_X1 _28948_ (.A(_05746_),
    .B1(_05889_),
    .B2(_05892_),
    .ZN(_05893_));
 NAND2_X1 _28949_ (.A1(_05738_),
    .A2(_05773_),
    .ZN(_05894_));
 AOI221_X2 _28950_ (.A(_05646_),
    .B1(_05821_),
    .B2(_05642_),
    .C1(_05894_),
    .C2(_05623_),
    .ZN(_05895_));
 OR3_X1 _28951_ (.A1(_05746_),
    .A2(_05672_),
    .A3(_05895_),
    .ZN(_05896_));
 AND4_X1 _28952_ (.A1(_05650_),
    .A2(_05886_),
    .A3(_05893_),
    .A4(_05896_),
    .ZN(_05897_));
 NAND2_X1 _28953_ (.A1(_05778_),
    .A2(_05767_),
    .ZN(_05898_));
 NOR2_X1 _28954_ (.A1(_15315_),
    .A2(_05898_),
    .ZN(_05899_));
 AND2_X1 _28955_ (.A1(_05728_),
    .A2(_05734_),
    .ZN(_05900_));
 NOR3_X1 _28956_ (.A1(_15308_),
    .A2(_05900_),
    .A3(_05774_),
    .ZN(_05901_));
 OAI21_X1 _28957_ (.A(_05640_),
    .B1(_05899_),
    .B2(_05901_),
    .ZN(_05902_));
 NAND3_X1 _28958_ (.A1(_05759_),
    .A2(_05750_),
    .A3(_05773_),
    .ZN(_05903_));
 AOI21_X4 _28959_ (.A(_05727_),
    .B1(_05598_),
    .B2(_05603_),
    .ZN(_05904_));
 OAI21_X1 _28960_ (.A(_15308_),
    .B1(_05872_),
    .B2(_05904_),
    .ZN(_05905_));
 NAND3_X1 _28961_ (.A1(_05715_),
    .A2(_05903_),
    .A3(_05905_),
    .ZN(_05906_));
 AOI21_X1 _28962_ (.A(_05714_),
    .B1(_05759_),
    .B2(_05841_),
    .ZN(_05907_));
 AOI21_X1 _28963_ (.A(_05904_),
    .B1(_05696_),
    .B2(_05704_),
    .ZN(_05908_));
 OAI21_X1 _28964_ (.A(_05907_),
    .B1(_05908_),
    .B2(_15315_),
    .ZN(_05909_));
 NAND3_X1 _28965_ (.A1(_05650_),
    .A2(_05906_),
    .A3(_05909_),
    .ZN(_05910_));
 NOR2_X1 _28966_ (.A1(_05639_),
    .A2(_05671_),
    .ZN(_05911_));
 AOI21_X4 _28967_ (.A(_05549_),
    .B1(_05598_),
    .B2(_05603_),
    .ZN(_05912_));
 NOR3_X4 _28968_ (.A1(_05727_),
    .A2(_05656_),
    .A3(_05657_),
    .ZN(_05913_));
 NOR3_X1 _28969_ (.A1(_05759_),
    .A2(_05912_),
    .A3(_05913_),
    .ZN(_05914_));
 AOI21_X4 _28970_ (.A(net1028),
    .B1(_05598_),
    .B2(_05603_),
    .ZN(_05915_));
 AOI21_X1 _28971_ (.A(_05915_),
    .B1(_05701_),
    .B2(_15296_),
    .ZN(_05916_));
 AOI21_X1 _28972_ (.A(_05914_),
    .B1(_05916_),
    .B2(_15315_),
    .ZN(_05917_));
 NAND2_X1 _28973_ (.A1(_05911_),
    .A2(_05917_),
    .ZN(_05918_));
 NAND3_X1 _28974_ (.A1(_05902_),
    .A2(_05910_),
    .A3(_05918_),
    .ZN(_05919_));
 OAI222_X2 _28975_ (.A1(_05851_),
    .A2(_05866_),
    .B1(_05882_),
    .B2(_05897_),
    .C1(_05919_),
    .C2(_05582_),
    .ZN(_00154_));
 NAND2_X2 _28976_ (.A1(_05549_),
    .A2(_05563_),
    .ZN(_05920_));
 AOI221_X2 _28977_ (.A(_05670_),
    .B1(_05598_),
    .B2(_05603_),
    .C1(_05564_),
    .C2(net101),
    .ZN(_05921_));
 NAND2_X1 _28978_ (.A1(_05727_),
    .A2(_05623_),
    .ZN(_05922_));
 OAI21_X1 _28979_ (.A(_05922_),
    .B1(_05876_),
    .B2(_05623_),
    .ZN(_05923_));
 NAND2_X1 _28980_ (.A1(_05632_),
    .A2(_05923_),
    .ZN(_05924_));
 NOR2_X1 _28981_ (.A1(_05591_),
    .A2(_05846_),
    .ZN(_05925_));
 AOI221_X2 _28982_ (.A(_05621_),
    .B1(_05920_),
    .B2(_05921_),
    .C1(_05924_),
    .C2(_05925_),
    .ZN(_05926_));
 OAI21_X1 _28983_ (.A(_05570_),
    .B1(_05757_),
    .B2(_05913_),
    .ZN(_05927_));
 OAI21_X1 _28984_ (.A(_05740_),
    .B1(_05754_),
    .B2(_05915_),
    .ZN(_05928_));
 NAND3_X1 _28985_ (.A1(_05911_),
    .A2(_05927_),
    .A3(_05928_),
    .ZN(_05929_));
 OAI21_X1 _28986_ (.A(_05568_),
    .B1(_05631_),
    .B2(_05532_),
    .ZN(_05930_));
 AOI221_X2 _28987_ (.A(_05737_),
    .B1(_05930_),
    .B2(_05549_),
    .C1(_05723_),
    .C2(_05533_),
    .ZN(_05931_));
 OAI21_X1 _28988_ (.A(_05929_),
    .B1(_05931_),
    .B2(_05782_),
    .ZN(_05932_));
 AOI221_X2 _28989_ (.A(_05591_),
    .B1(_05920_),
    .B2(_05729_),
    .C1(_05631_),
    .C2(_05568_),
    .ZN(_05933_));
 NOR3_X1 _28990_ (.A1(_05568_),
    .A2(_05666_),
    .A3(_05904_),
    .ZN(_05934_));
 AOI21_X2 _28991_ (.A(_05867_),
    .B1(_05631_),
    .B2(_05531_),
    .ZN(_05935_));
 AOI21_X2 _28992_ (.A(_05934_),
    .B1(_05935_),
    .B2(_05569_),
    .ZN(_05936_));
 AOI211_X2 _28993_ (.A(_05621_),
    .B(_05933_),
    .C1(_05936_),
    .C2(_05713_),
    .ZN(_05937_));
 AOI22_X1 _28994_ (.A1(_05719_),
    .A2(_05592_),
    .B1(_05679_),
    .B2(_05567_),
    .ZN(_05938_));
 OAI221_X1 _28995_ (.A(_05640_),
    .B1(_05938_),
    .B2(_05709_),
    .C1(_05644_),
    .C2(_05684_),
    .ZN(_05939_));
 AOI21_X1 _28996_ (.A(_05939_),
    .B1(_05724_),
    .B2(_05698_),
    .ZN(_05940_));
 NAND2_X1 _28997_ (.A1(_05683_),
    .A2(_05724_),
    .ZN(_05941_));
 NAND2_X1 _28998_ (.A1(net103),
    .A2(_05872_),
    .ZN(_05942_));
 NAND4_X2 _28999_ (.A1(_05911_),
    .A2(_05868_),
    .A3(_05941_),
    .A4(_05942_),
    .ZN(_05943_));
 NAND3_X2 _29000_ (.A1(_05943_),
    .A2(_05581_),
    .A3(_05676_),
    .ZN(_05944_));
 OAI33_X1 _29001_ (.A1(_05582_),
    .A2(_05926_),
    .A3(_05932_),
    .B1(_05937_),
    .B2(_05940_),
    .B3(_05944_),
    .ZN(_05945_));
 NOR2_X1 _29002_ (.A1(_05676_),
    .A2(_05746_),
    .ZN(_05946_));
 AOI22_X1 _29003_ (.A1(_05755_),
    .A2(_05703_),
    .B1(_05822_),
    .B2(_05728_),
    .ZN(_05947_));
 OAI21_X1 _29004_ (.A(_05946_),
    .B1(_05947_),
    .B2(_05782_),
    .ZN(_05948_));
 INV_X1 _29005_ (.A(_05948_),
    .ZN(_05949_));
 AOI21_X1 _29006_ (.A(_05569_),
    .B1(_05655_),
    .B2(_05778_),
    .ZN(_05950_));
 AOI21_X1 _29007_ (.A(_05757_),
    .B1(_05876_),
    .B2(_05632_),
    .ZN(_05951_));
 AOI21_X1 _29008_ (.A(_05950_),
    .B1(_05951_),
    .B2(_05570_),
    .ZN(_05952_));
 NOR3_X1 _29009_ (.A1(_05733_),
    .A2(_05718_),
    .A3(_05952_),
    .ZN(_05953_));
 OAI21_X1 _29010_ (.A(_05621_),
    .B1(_05656_),
    .B2(_05657_),
    .ZN(_05954_));
 OAI22_X1 _29011_ (.A1(_05740_),
    .A2(_05954_),
    .B1(_05702_),
    .B2(_05734_),
    .ZN(_05955_));
 NOR2_X1 _29012_ (.A1(_05696_),
    .A2(_05702_),
    .ZN(_05956_));
 AOI22_X1 _29013_ (.A1(_05698_),
    .A2(_05955_),
    .B1(_05956_),
    .B2(_05684_),
    .ZN(_05957_));
 NAND2_X1 _29014_ (.A1(_05634_),
    .A2(_05696_),
    .ZN(_05958_));
 NAND3_X1 _29015_ (.A1(net103),
    .A2(_05639_),
    .A3(_05720_),
    .ZN(_05959_));
 AND2_X1 _29016_ (.A1(_05958_),
    .A2(_05959_),
    .ZN(_05960_));
 OAI21_X1 _29017_ (.A(_05957_),
    .B1(_05960_),
    .B2(_05759_),
    .ZN(_05961_));
 AOI21_X2 _29018_ (.A(_05953_),
    .B1(_05961_),
    .B2(_05715_),
    .ZN(_05962_));
 NOR3_X1 _29019_ (.A1(_15296_),
    .A2(_05717_),
    .A3(_05703_),
    .ZN(_05963_));
 AOI21_X1 _29020_ (.A(_05625_),
    .B1(_05883_),
    .B2(_15290_),
    .ZN(_05964_));
 OAI21_X1 _29021_ (.A(_05755_),
    .B1(_05963_),
    .B2(_05964_),
    .ZN(_05965_));
 NAND2_X1 _29022_ (.A1(_05740_),
    .A2(_05883_),
    .ZN(_05966_));
 XNOR2_X1 _29023_ (.A(_05633_),
    .B(_05713_),
    .ZN(_05967_));
 OAI221_X1 _29024_ (.A(_05701_),
    .B1(_05966_),
    .B2(_15296_),
    .C1(_05967_),
    .C2(net902),
    .ZN(_05968_));
 NAND3_X1 _29025_ (.A1(_15299_),
    .A2(_15308_),
    .A3(_05718_),
    .ZN(_05969_));
 NAND4_X1 _29026_ (.A1(_05649_),
    .A2(_05965_),
    .A3(_05968_),
    .A4(_05969_),
    .ZN(_05970_));
 AOI21_X1 _29027_ (.A(_05789_),
    .B1(_05748_),
    .B2(_05683_),
    .ZN(_05971_));
 OR2_X1 _29028_ (.A1(_05661_),
    .A2(_05774_),
    .ZN(_05972_));
 MUX2_X1 _29029_ (.A(_05971_),
    .B(_05972_),
    .S(_05566_),
    .Z(_05973_));
 NOR3_X1 _29030_ (.A1(_05566_),
    .A2(_05666_),
    .A3(_05867_),
    .ZN(_05974_));
 AOI21_X1 _29031_ (.A(_05665_),
    .B1(_05658_),
    .B2(_05750_),
    .ZN(_05975_));
 OR2_X1 _29032_ (.A1(_05974_),
    .A2(_05975_),
    .ZN(_05976_));
 OAI221_X2 _29033_ (.A(_05970_),
    .B1(_05973_),
    .B2(_05787_),
    .C1(_05782_),
    .C2(_05976_),
    .ZN(_05977_));
 AND2_X1 _29034_ (.A1(_05575_),
    .A2(_05581_),
    .ZN(_05978_));
 AOI221_X2 _29035_ (.A(_05945_),
    .B1(_05949_),
    .B2(_05962_),
    .C1(_05977_),
    .C2(_05978_),
    .ZN(_00155_));
 NOR3_X2 _29036_ (.A1(_05757_),
    .A2(_05633_),
    .A3(_05913_),
    .ZN(_05979_));
 NOR2_X1 _29037_ (.A1(_05740_),
    .A2(_05915_),
    .ZN(_05980_));
 NAND2_X4 _29038_ (.A1(_05533_),
    .A2(_05872_),
    .ZN(_05981_));
 AOI21_X1 _29039_ (.A(_05979_),
    .B1(_05980_),
    .B2(_05981_),
    .ZN(_05982_));
 AND2_X1 _29040_ (.A1(_05727_),
    .A2(_05633_),
    .ZN(_05983_));
 AOI21_X1 _29041_ (.A(_05983_),
    .B1(_05825_),
    .B2(_05566_),
    .ZN(_05984_));
 OAI221_X1 _29042_ (.A(_05978_),
    .B1(_05982_),
    .B2(_05782_),
    .C1(_05984_),
    .C2(_05787_),
    .ZN(_05985_));
 NOR2_X1 _29043_ (.A1(_05623_),
    .A2(_05765_),
    .ZN(_05986_));
 AOI21_X2 _29044_ (.A(_05915_),
    .B1(_05631_),
    .B2(net100),
    .ZN(_05987_));
 AOI221_X2 _29045_ (.A(_05671_),
    .B1(_05986_),
    .B2(_05981_),
    .C1(_05987_),
    .C2(_05624_),
    .ZN(_05988_));
 OAI21_X1 _29046_ (.A(_05625_),
    .B1(_05566_),
    .B2(_15292_),
    .ZN(_05989_));
 NAND2_X1 _29047_ (.A1(_05701_),
    .A2(_05989_),
    .ZN(_05990_));
 AOI21_X2 _29048_ (.A(_05988_),
    .B1(_05990_),
    .B2(_05736_),
    .ZN(_05991_));
 AOI21_X2 _29049_ (.A(_05985_),
    .B1(_05991_),
    .B2(_05650_),
    .ZN(_05992_));
 NOR2_X1 _29050_ (.A1(net910),
    .A2(_05620_),
    .ZN(_05993_));
 AOI221_X2 _29051_ (.A(_05670_),
    .B1(_05662_),
    .B2(_05993_),
    .C1(_05912_),
    .C2(_05533_),
    .ZN(_05994_));
 AOI21_X1 _29052_ (.A(_05913_),
    .B1(_05720_),
    .B2(_05622_),
    .ZN(_05995_));
 OAI21_X1 _29053_ (.A(_05994_),
    .B1(_05995_),
    .B2(_05802_),
    .ZN(_05996_));
 OAI21_X1 _29054_ (.A(_05692_),
    .B1(_05644_),
    .B2(_05693_),
    .ZN(_05997_));
 AOI21_X1 _29055_ (.A(_05996_),
    .B1(_05997_),
    .B2(net105),
    .ZN(_05998_));
 NOR2_X1 _29056_ (.A1(_05677_),
    .A2(_05998_),
    .ZN(_05999_));
 MUX2_X1 _29057_ (.A(_15304_),
    .B(_05817_),
    .S(_05696_),
    .Z(_06000_));
 NAND2_X1 _29058_ (.A1(_05733_),
    .A2(_06000_),
    .ZN(_06001_));
 OAI21_X1 _29059_ (.A(_05981_),
    .B1(_05680_),
    .B2(_05634_),
    .ZN(_06002_));
 AOI21_X1 _29060_ (.A(_05665_),
    .B1(_05738_),
    .B2(_05783_),
    .ZN(_06003_));
 OAI21_X1 _29061_ (.A(_05649_),
    .B1(_06002_),
    .B2(_06003_),
    .ZN(_06004_));
 NAND3_X1 _29062_ (.A1(_05673_),
    .A2(_06001_),
    .A3(_06004_),
    .ZN(_06005_));
 NOR3_X1 _29063_ (.A1(net100),
    .A2(_05623_),
    .A3(_05591_),
    .ZN(_06006_));
 NOR2_X1 _29064_ (.A1(_05568_),
    .A2(_05670_),
    .ZN(_06007_));
 AOI21_X1 _29065_ (.A(_06006_),
    .B1(_06007_),
    .B2(_15292_),
    .ZN(_06008_));
 OAI21_X1 _29066_ (.A(net910),
    .B1(_05568_),
    .B2(_05591_),
    .ZN(_06009_));
 AOI21_X1 _29067_ (.A(_05592_),
    .B1(_06009_),
    .B2(_05533_),
    .ZN(_06010_));
 MUX2_X1 _29068_ (.A(_06008_),
    .B(_06010_),
    .S(_05719_),
    .Z(_06011_));
 OAI22_X1 _29069_ (.A1(_05624_),
    .A2(_05671_),
    .B1(_05719_),
    .B2(_05763_),
    .ZN(_06012_));
 AOI21_X1 _29070_ (.A(_05814_),
    .B1(_06012_),
    .B2(_05704_),
    .ZN(_06013_));
 NOR2_X1 _29071_ (.A1(_05663_),
    .A2(_05563_),
    .ZN(_06014_));
 OAI21_X1 _29072_ (.A(_05734_),
    .B1(_05842_),
    .B2(_06014_),
    .ZN(_06015_));
 AOI22_X2 _29073_ (.A1(_05776_),
    .A2(_06007_),
    .B1(_06015_),
    .B2(_05607_),
    .ZN(_06016_));
 NOR2_X2 _29074_ (.A1(_05581_),
    .A2(_05693_),
    .ZN(_06017_));
 AOI221_X2 _29075_ (.A(_05576_),
    .B1(_06011_),
    .B2(_06013_),
    .C1(_06016_),
    .C2(_06017_),
    .ZN(_06018_));
 AOI21_X1 _29076_ (.A(_05569_),
    .B1(_05631_),
    .B2(_05533_),
    .ZN(_06019_));
 AOI21_X1 _29077_ (.A(_05592_),
    .B1(_05783_),
    .B2(_06019_),
    .ZN(_06020_));
 AOI21_X1 _29078_ (.A(_05671_),
    .B1(_05696_),
    .B2(_05728_),
    .ZN(_06021_));
 AOI221_X2 _29079_ (.A(_05828_),
    .B1(_06020_),
    .B2(_05883_),
    .C1(_06021_),
    .C2(_05790_),
    .ZN(_06022_));
 OAI21_X1 _29080_ (.A(_05750_),
    .B1(_05632_),
    .B2(_15292_),
    .ZN(_06023_));
 XNOR2_X1 _29081_ (.A(_05533_),
    .B(_05631_),
    .ZN(_06024_));
 MUX2_X1 _29082_ (.A(_06023_),
    .B(_06024_),
    .S(_05624_),
    .Z(_06025_));
 OAI22_X1 _29083_ (.A1(_15299_),
    .A2(_05680_),
    .B1(_05915_),
    .B2(_05570_),
    .ZN(_06026_));
 MUX2_X1 _29084_ (.A(_06025_),
    .B(_06026_),
    .S(_05672_),
    .Z(_06027_));
 NOR2_X1 _29085_ (.A1(_05581_),
    .A2(_05622_),
    .ZN(_06028_));
 AOI21_X2 _29086_ (.A(_06022_),
    .B1(_06027_),
    .B2(_06028_),
    .ZN(_06029_));
 AOI221_X2 _29087_ (.A(_05992_),
    .B1(_05999_),
    .B2(_06005_),
    .C1(_06018_),
    .C2(_06029_),
    .ZN(_00156_));
 NOR2_X1 _29088_ (.A1(_05633_),
    .A2(_05904_),
    .ZN(_06030_));
 AOI21_X1 _29089_ (.A(_05774_),
    .B1(_05748_),
    .B2(_05704_),
    .ZN(_06031_));
 AOI221_X2 _29090_ (.A(_05883_),
    .B1(_05981_),
    .B2(_06030_),
    .C1(_06031_),
    .C2(_05802_),
    .ZN(_06032_));
 AOI221_X1 _29091_ (.A(_05714_),
    .B1(_05680_),
    .B2(_05549_),
    .C1(_05912_),
    .C2(_15296_),
    .ZN(_06033_));
 NOR3_X1 _29092_ (.A1(_05576_),
    .A2(_06032_),
    .A3(_06033_),
    .ZN(_06034_));
 NOR2_X1 _29093_ (.A1(_05605_),
    .A2(_05703_),
    .ZN(_06035_));
 OAI221_X1 _29094_ (.A(_05673_),
    .B1(_05644_),
    .B2(_05877_),
    .C1(_06035_),
    .C2(_05658_),
    .ZN(_06036_));
 NAND2_X1 _29095_ (.A1(_05642_),
    .A2(_05565_),
    .ZN(_06037_));
 AOI21_X1 _29096_ (.A(_05672_),
    .B1(_05755_),
    .B2(_06037_),
    .ZN(_06038_));
 OAI21_X1 _29097_ (.A(_06038_),
    .B1(_05810_),
    .B2(net101),
    .ZN(_06039_));
 AOI21_X1 _29098_ (.A(_05676_),
    .B1(_06036_),
    .B2(_06039_),
    .ZN(_06040_));
 OAI21_X1 _29099_ (.A(_06017_),
    .B1(_06034_),
    .B2(_06040_),
    .ZN(_06041_));
 AOI22_X2 _29100_ (.A1(_05734_),
    .A2(_05690_),
    .B1(_05692_),
    .B2(net103),
    .ZN(_06042_));
 AOI221_X2 _29101_ (.A(_05671_),
    .B1(_05679_),
    .B2(_05683_),
    .C1(_05821_),
    .C2(net910),
    .ZN(_06043_));
 NOR2_X1 _29102_ (.A1(net103),
    .A2(_05644_),
    .ZN(_06044_));
 OAI21_X1 _29103_ (.A(_15299_),
    .B1(_05651_),
    .B2(_06044_),
    .ZN(_06045_));
 AOI221_X2 _29104_ (.A(_05675_),
    .B1(_05883_),
    .B2(_06042_),
    .C1(_06043_),
    .C2(_06045_),
    .ZN(_06046_));
 OAI21_X1 _29105_ (.A(_05900_),
    .B1(_05729_),
    .B2(_05759_),
    .ZN(_06047_));
 NOR2_X1 _29106_ (.A1(_05576_),
    .A2(_05672_),
    .ZN(_06048_));
 AND4_X1 _29107_ (.A1(_05722_),
    .A2(_05750_),
    .A3(_06047_),
    .A4(_06048_),
    .ZN(_06049_));
 NAND2_X1 _29108_ (.A1(_05676_),
    .A2(_05673_),
    .ZN(_06050_));
 OAI21_X1 _29109_ (.A(_05658_),
    .B1(_05755_),
    .B2(net101),
    .ZN(_06051_));
 NOR2_X1 _29110_ (.A1(net654),
    .A2(_05748_),
    .ZN(_06052_));
 OAI22_X1 _29111_ (.A1(_15308_),
    .A2(_06051_),
    .B1(_06052_),
    .B2(_05790_),
    .ZN(_06053_));
 OAI21_X1 _29112_ (.A(_05799_),
    .B1(_06050_),
    .B2(_06053_),
    .ZN(_06054_));
 OR3_X1 _29113_ (.A1(_06046_),
    .A2(_06049_),
    .A3(_06054_),
    .ZN(_06055_));
 AOI22_X2 _29114_ (.A1(net654),
    .A2(_05755_),
    .B1(_05981_),
    .B2(_15315_),
    .ZN(_06056_));
 NAND2_X1 _29115_ (.A1(_05576_),
    .A2(_05581_),
    .ZN(_06057_));
 NOR3_X1 _29116_ (.A1(_05802_),
    .A2(_05789_),
    .A3(_05915_),
    .ZN(_06058_));
 NOR2_X2 _29117_ (.A1(_05664_),
    .A2(_05644_),
    .ZN(_06059_));
 NOR4_X2 _29118_ (.A1(_05715_),
    .A2(_06057_),
    .A3(_06058_),
    .A4(_06059_),
    .ZN(_06060_));
 AOI21_X1 _29119_ (.A(_05714_),
    .B1(_05679_),
    .B2(_15299_),
    .ZN(_06061_));
 AOI21_X1 _29120_ (.A(_05851_),
    .B1(_05927_),
    .B2(_06061_),
    .ZN(_06062_));
 OAI22_X2 _29121_ (.A1(_05673_),
    .A2(_06056_),
    .B1(_06060_),
    .B2(_06062_),
    .ZN(_06063_));
 AOI21_X1 _29122_ (.A(_05802_),
    .B1(_05749_),
    .B2(_05767_),
    .ZN(_06064_));
 NOR2_X1 _29123_ (.A1(_15296_),
    .A2(_05680_),
    .ZN(_06065_));
 OR3_X1 _29124_ (.A1(_06057_),
    .A2(_06064_),
    .A3(_06065_),
    .ZN(_06066_));
 AOI22_X1 _29125_ (.A1(_05683_),
    .A2(_05632_),
    .B1(_05690_),
    .B2(_05821_),
    .ZN(_06067_));
 NOR3_X1 _29126_ (.A1(_05675_),
    .A2(_05717_),
    .A3(_06067_),
    .ZN(_06068_));
 NOR4_X4 _29127_ (.A1(_05867_),
    .A2(_05675_),
    .A3(_05774_),
    .A4(_05564_),
    .ZN(_06069_));
 NOR2_X1 _29128_ (.A1(_05690_),
    .A2(_05680_),
    .ZN(_06070_));
 OAI21_X1 _29129_ (.A(_05773_),
    .B1(_05604_),
    .B2(_05683_),
    .ZN(_06071_));
 AOI221_X2 _29130_ (.A(_06069_),
    .B1(_06070_),
    .B2(_05675_),
    .C1(_06071_),
    .C2(_05565_),
    .ZN(_06072_));
 AOI21_X1 _29131_ (.A(_05696_),
    .B1(_05920_),
    .B2(_06037_),
    .ZN(_06073_));
 NOR2_X1 _29132_ (.A1(_05576_),
    .A2(_06073_),
    .ZN(_06074_));
 AOI221_X2 _29133_ (.A(_06068_),
    .B1(_06072_),
    .B2(_05714_),
    .C1(_05607_),
    .C2(_06074_),
    .ZN(_06075_));
 OAI221_X2 _29134_ (.A(_06063_),
    .B1(_06066_),
    .B2(_05673_),
    .C1(_06075_),
    .C2(_05746_),
    .ZN(_06076_));
 OAI211_X2 _29135_ (.A(_06041_),
    .B(_06055_),
    .C1(_06076_),
    .C2(_05733_),
    .ZN(_00157_));
 NAND2_X1 _29136_ (.A1(_05883_),
    .A2(_05867_),
    .ZN(_06077_));
 OAI21_X1 _29137_ (.A(_05696_),
    .B1(_05713_),
    .B2(_05728_),
    .ZN(_06078_));
 NAND3_X1 _29138_ (.A1(_05665_),
    .A2(_06077_),
    .A3(_06078_),
    .ZN(_06079_));
 OAI221_X2 _29139_ (.A(_05740_),
    .B1(_05720_),
    .B2(_05763_),
    .C1(_05883_),
    .C2(_05534_),
    .ZN(_06080_));
 AOI221_X2 _29140_ (.A(_05622_),
    .B1(_05714_),
    .B2(_05661_),
    .C1(_06079_),
    .C2(_06080_),
    .ZN(_06081_));
 NOR3_X1 _29141_ (.A1(_05709_),
    .A2(_05549_),
    .A3(_05591_),
    .ZN(_06082_));
 OR2_X2 _29142_ (.A1(_05670_),
    .A2(_05915_),
    .ZN(_06083_));
 NOR2_X1 _29143_ (.A1(_05713_),
    .A2(_05734_),
    .ZN(_06084_));
 AOI221_X2 _29144_ (.A(_06082_),
    .B1(_06083_),
    .B2(_05857_),
    .C1(_05703_),
    .C2(_06084_),
    .ZN(_06085_));
 NOR4_X1 _29145_ (.A1(_05527_),
    .A2(_05530_),
    .A3(_05549_),
    .A4(_05565_),
    .ZN(_06086_));
 OAI21_X1 _29146_ (.A(_05818_),
    .B1(_05661_),
    .B2(_06086_),
    .ZN(_06087_));
 AND3_X1 _29147_ (.A1(_05710_),
    .A2(_05942_),
    .A3(_06087_),
    .ZN(_06088_));
 OAI22_X1 _29148_ (.A1(_05650_),
    .A2(_06085_),
    .B1(_06088_),
    .B2(_05787_),
    .ZN(_06089_));
 NOR3_X1 _29149_ (.A1(_05582_),
    .A2(_06081_),
    .A3(_06089_),
    .ZN(_06090_));
 AOI21_X1 _29150_ (.A(_05913_),
    .B1(_05720_),
    .B2(_05683_),
    .ZN(_06091_));
 OAI221_X1 _29151_ (.A(_05714_),
    .B1(_05644_),
    .B2(_05534_),
    .C1(_06091_),
    .C2(_05665_),
    .ZN(_06092_));
 AND3_X1 _29152_ (.A1(_05649_),
    .A2(_05884_),
    .A3(_06092_),
    .ZN(_06093_));
 NAND2_X1 _29153_ (.A1(_15310_),
    .A2(_05742_),
    .ZN(_06094_));
 OAI221_X2 _29154_ (.A(_05922_),
    .B1(_05657_),
    .B2(_05656_),
    .C1(_05704_),
    .C2(_05740_),
    .ZN(_06095_));
 AOI21_X1 _29155_ (.A(_05782_),
    .B1(_06094_),
    .B2(_06095_),
    .ZN(_06096_));
 NOR3_X1 _29156_ (.A1(_05787_),
    .A2(_05950_),
    .A3(_06059_),
    .ZN(_06097_));
 OR2_X1 _29157_ (.A1(_06096_),
    .A2(_06097_),
    .ZN(_06098_));
 NOR3_X1 _29158_ (.A1(_05867_),
    .A2(_05754_),
    .A3(_05665_),
    .ZN(_06099_));
 AOI221_X2 _29159_ (.A(_05565_),
    .B1(_05604_),
    .B2(_05876_),
    .C1(_05872_),
    .C2(_05533_),
    .ZN(_06100_));
 NOR4_X2 _29160_ (.A1(_06099_),
    .A2(_05718_),
    .A3(_06100_),
    .A4(_05733_),
    .ZN(_06101_));
 NOR2_X1 _29161_ (.A1(_15294_),
    .A2(_05631_),
    .ZN(_06102_));
 NOR2_X1 _29162_ (.A1(_05569_),
    .A2(_06102_),
    .ZN(_06103_));
 AOI221_X2 _29163_ (.A(_05782_),
    .B1(_05981_),
    .B2(_06103_),
    .C1(_05935_),
    .C2(_05570_),
    .ZN(_06104_));
 OAI221_X1 _29164_ (.A(_05734_),
    .B1(_05645_),
    .B2(_05709_),
    .C1(_05624_),
    .C2(net102),
    .ZN(_06105_));
 OAI21_X1 _29165_ (.A(_06105_),
    .B1(_05748_),
    .B2(_15311_),
    .ZN(_06106_));
 OAI21_X1 _29166_ (.A(_05696_),
    .B1(_05703_),
    .B2(_05704_),
    .ZN(_06107_));
 NAND2_X1 _29167_ (.A1(_05725_),
    .A2(_06107_),
    .ZN(_06108_));
 OAI221_X1 _29168_ (.A(_05978_),
    .B1(_06106_),
    .B2(_05787_),
    .C1(_06108_),
    .C2(_05840_),
    .ZN(_06109_));
 OAI33_X1 _29169_ (.A1(_05677_),
    .A2(_06093_),
    .A3(_06098_),
    .B1(_06101_),
    .B2(_06104_),
    .B3(_06109_),
    .ZN(_06110_));
 AOI21_X1 _29170_ (.A(_05759_),
    .B1(_05958_),
    .B2(_05773_),
    .ZN(_06111_));
 OAI22_X1 _29171_ (.A1(_05728_),
    .A2(_05742_),
    .B1(_05738_),
    .B2(_05704_),
    .ZN(_06112_));
 OAI21_X1 _29172_ (.A(_05672_),
    .B1(_06112_),
    .B2(_05802_),
    .ZN(_06113_));
 AOI21_X2 _29173_ (.A(_05912_),
    .B1(_05742_),
    .B2(_05728_),
    .ZN(_06114_));
 NOR2_X1 _29174_ (.A1(_15315_),
    .A2(_06114_),
    .ZN(_06115_));
 OAI21_X1 _29175_ (.A(_05718_),
    .B1(_05810_),
    .B2(_05841_),
    .ZN(_06116_));
 OAI221_X1 _29176_ (.A(_05650_),
    .B1(_06111_),
    .B2(_06113_),
    .C1(_06115_),
    .C2(_06116_),
    .ZN(_06117_));
 NAND2_X1 _29177_ (.A1(_05802_),
    .A2(_05733_),
    .ZN(_06118_));
 OAI21_X1 _29178_ (.A(_05783_),
    .B1(_05748_),
    .B2(_05728_),
    .ZN(_06119_));
 AOI22_X1 _29179_ (.A1(_05634_),
    .A2(_05742_),
    .B1(_05757_),
    .B2(_05693_),
    .ZN(_06120_));
 OAI22_X1 _29180_ (.A1(_06118_),
    .A2(_06119_),
    .B1(_06120_),
    .B2(_15308_),
    .ZN(_06121_));
 NOR2_X1 _29181_ (.A1(_05534_),
    .A2(_05740_),
    .ZN(_06122_));
 OR2_X1 _29182_ (.A1(_05794_),
    .A2(_06122_),
    .ZN(_06123_));
 NOR3_X1 _29183_ (.A1(_15309_),
    .A2(_15318_),
    .A3(_05742_),
    .ZN(_06124_));
 NOR2_X1 _29184_ (.A1(_05782_),
    .A2(_06124_),
    .ZN(_06125_));
 AOI22_X1 _29185_ (.A1(_05715_),
    .A2(_06121_),
    .B1(_06123_),
    .B2(_06125_),
    .ZN(_06126_));
 AOI21_X1 _29186_ (.A(_05851_),
    .B1(_06117_),
    .B2(_06126_),
    .ZN(_06127_));
 OR3_X2 _29187_ (.A1(_06110_),
    .A2(_06090_),
    .A3(_06127_),
    .ZN(_00158_));
 AOI221_X1 _29188_ (.A(_05883_),
    .B1(_05662_),
    .B2(_15292_),
    .C1(_05724_),
    .C2(_15290_),
    .ZN(_06128_));
 AOI21_X1 _29189_ (.A(_05912_),
    .B1(_05679_),
    .B2(_15299_),
    .ZN(_06129_));
 OAI21_X1 _29190_ (.A(_06128_),
    .B1(_06129_),
    .B2(net105),
    .ZN(_06130_));
 OAI221_X1 _29191_ (.A(_05673_),
    .B1(_05810_),
    .B2(_05728_),
    .C1(_05987_),
    .C2(_15315_),
    .ZN(_06131_));
 AND3_X1 _29192_ (.A1(_05747_),
    .A2(_06130_),
    .A3(_06131_),
    .ZN(_06132_));
 OAI222_X2 _29193_ (.A1(net101),
    .A2(_05644_),
    .B1(_05692_),
    .B2(_15299_),
    .C1(_05822_),
    .C2(_05664_),
    .ZN(_06133_));
 NAND3_X1 _29194_ (.A1(_05665_),
    .A2(_05738_),
    .A3(_05773_),
    .ZN(_06134_));
 OAI21_X1 _29195_ (.A(_06134_),
    .B1(_05908_),
    .B2(_05802_),
    .ZN(_06135_));
 MUX2_X1 _29196_ (.A(_06133_),
    .B(_06135_),
    .S(_05672_),
    .Z(_06136_));
 AND2_X1 _29197_ (.A1(_05762_),
    .A2(_06136_),
    .ZN(_06137_));
 NAND2_X1 _29198_ (.A1(_15296_),
    .A2(_05912_),
    .ZN(_06138_));
 OAI21_X1 _29199_ (.A(net105),
    .B1(_05724_),
    .B2(_05754_),
    .ZN(_06139_));
 AOI21_X1 _29200_ (.A(_05718_),
    .B1(_06138_),
    .B2(_06139_),
    .ZN(_06140_));
 AOI21_X1 _29201_ (.A(_05679_),
    .B1(_05703_),
    .B2(_05748_),
    .ZN(_06141_));
 AOI21_X1 _29202_ (.A(_05661_),
    .B1(_05662_),
    .B2(_15290_),
    .ZN(_06142_));
 OAI22_X1 _29203_ (.A1(net105),
    .A2(_06141_),
    .B1(_06142_),
    .B2(_05672_),
    .ZN(_06143_));
 OAI21_X1 _29204_ (.A(_06017_),
    .B1(_06140_),
    .B2(_06143_),
    .ZN(_06144_));
 AND2_X1 _29205_ (.A1(_05966_),
    .A2(_06028_),
    .ZN(_06145_));
 NOR3_X1 _29206_ (.A1(_05549_),
    .A2(_05671_),
    .A3(_05644_),
    .ZN(_06146_));
 OAI21_X1 _29207_ (.A(_05692_),
    .B1(_05720_),
    .B2(_05717_),
    .ZN(_06147_));
 AOI21_X1 _29208_ (.A(_06146_),
    .B1(_06147_),
    .B2(_15299_),
    .ZN(_06148_));
 OAI221_X1 _29209_ (.A(_06145_),
    .B1(_06148_),
    .B2(net105),
    .C1(_05698_),
    .C2(_05680_),
    .ZN(_06149_));
 AND3_X1 _29210_ (.A1(_05582_),
    .A2(_06144_),
    .A3(_06149_),
    .ZN(_06150_));
 NOR2_X1 _29211_ (.A1(_15318_),
    .A2(_05720_),
    .ZN(_06151_));
 AOI221_X1 _29212_ (.A(_06014_),
    .B1(_05654_),
    .B2(_05653_),
    .C1(_05727_),
    .C2(_05569_),
    .ZN(_06152_));
 OAI21_X1 _29213_ (.A(_05693_),
    .B1(_06151_),
    .B2(_06152_),
    .ZN(_06153_));
 NAND2_X1 _29214_ (.A1(_05634_),
    .A2(_05623_),
    .ZN(_06154_));
 MUX2_X1 _29215_ (.A(_15304_),
    .B(_06154_),
    .S(_05719_),
    .Z(_06155_));
 AOI21_X1 _29216_ (.A(_05717_),
    .B1(_06155_),
    .B2(_05622_),
    .ZN(_06156_));
 MUX2_X1 _29217_ (.A(_05698_),
    .B(_05642_),
    .S(_05620_),
    .Z(_06157_));
 OAI33_X1 _29218_ (.A1(_05693_),
    .A2(_05658_),
    .A3(_05703_),
    .B1(_06157_),
    .B2(_05734_),
    .B3(_05624_),
    .ZN(_06158_));
 OAI21_X1 _29219_ (.A(_05714_),
    .B1(_05702_),
    .B2(_05898_),
    .ZN(_06159_));
 NOR2_X1 _29220_ (.A1(_06158_),
    .A2(_06159_),
    .ZN(_06160_));
 MUX2_X1 _29221_ (.A(_05679_),
    .B(_05821_),
    .S(_05639_),
    .Z(_06161_));
 NAND2_X1 _29222_ (.A1(net105),
    .A2(_06161_),
    .ZN(_06162_));
 AOI221_X2 _29223_ (.A(_05676_),
    .B1(_06153_),
    .B2(_06156_),
    .C1(_06160_),
    .C2(_06162_),
    .ZN(_06163_));
 OAI221_X1 _29224_ (.A(_05830_),
    .B1(_05644_),
    .B2(_05876_),
    .C1(_06114_),
    .C2(_05802_),
    .ZN(_06164_));
 AND2_X1 _29225_ (.A1(_05733_),
    .A2(_06164_),
    .ZN(_06165_));
 OAI221_X1 _29226_ (.A(_05649_),
    .B1(_05794_),
    .B2(_06122_),
    .C1(_05701_),
    .C2(net654),
    .ZN(_06166_));
 NAND2_X1 _29227_ (.A1(_06048_),
    .A2(_06166_),
    .ZN(_06167_));
 OAI21_X1 _29228_ (.A(_05746_),
    .B1(_06165_),
    .B2(_06167_),
    .ZN(_06168_));
 NAND3_X1 _29229_ (.A1(_05566_),
    .A2(_05694_),
    .A3(_05803_),
    .ZN(_06169_));
 NAND3_X1 _29230_ (.A1(_05733_),
    .A2(_05806_),
    .A3(_06169_),
    .ZN(_06170_));
 OAI21_X1 _29231_ (.A(_05624_),
    .B1(_05734_),
    .B2(_05709_),
    .ZN(_06171_));
 OAI221_X2 _29232_ (.A(_05693_),
    .B1(_06102_),
    .B2(_06171_),
    .C1(_05566_),
    .C2(_15292_),
    .ZN(_06172_));
 AOI221_X1 _29233_ (.A(_05576_),
    .B1(_05585_),
    .B2(_05589_),
    .C1(_06170_),
    .C2(_06172_),
    .ZN(_06173_));
 OAI33_X1 _29234_ (.A1(_06132_),
    .A2(_06137_),
    .A3(_06150_),
    .B1(_06163_),
    .B2(_06168_),
    .B3(_06173_),
    .ZN(_00159_));
 BUF_X1 _29235_ (.A(\dcnt[0] ),
    .Z(_06174_));
 BUF_X1 _29236_ (.A(\dcnt[2] ),
    .Z(_06175_));
 NOR3_X1 _29237_ (.A1(\dcnt[1] ),
    .A2(\dcnt[3] ),
    .A3(_06175_),
    .ZN(_06176_));
 AND3_X1 _29238_ (.A1(_06797_),
    .A2(_06174_),
    .A3(_06176_),
    .ZN(_00160_));
 XOR2_X2 _29239_ (.A(_06598_),
    .B(\sa00_sr[0] ),
    .Z(_00185_));
 XOR2_X2 _29240_ (.A(_06614_),
    .B(net839),
    .Z(_00186_));
 XOR2_X2 _29241_ (.A(_06630_),
    .B(_09088_),
    .Z(_00187_));
 XOR2_X2 _29242_ (.A(_06649_),
    .B(_09186_),
    .Z(_00188_));
 XOR2_X2 _29243_ (.A(_06666_),
    .B(_09162_),
    .Z(_00189_));
 XOR2_X2 _29244_ (.A(_06683_),
    .B(_09065_),
    .Z(_00190_));
 XOR2_X2 _29245_ (.A(_06701_),
    .B(_09154_),
    .Z(_00191_));
 XOR2_X1 _29246_ (.A(_06706_),
    .B(_08978_),
    .Z(_00192_));
 XOR2_X1 _29247_ (.A(net784),
    .B(_09719_),
    .Z(_00281_));
 XOR2_X1 _29248_ (.A(net1089),
    .B(net753),
    .Z(_00282_));
 XOR2_X1 _29249_ (.A(_06638_),
    .B(_09835_),
    .Z(_00283_));
 XOR2_X1 _29250_ (.A(_06657_),
    .B(_09868_),
    .Z(_00284_));
 XOR2_X1 _29251_ (.A(_06673_),
    .B(_09813_),
    .Z(_00285_));
 XOR2_X1 _29252_ (.A(_06688_),
    .B(_09789_),
    .Z(_00286_));
 XOR2_X1 _29253_ (.A(_06697_),
    .B(_09798_),
    .Z(_00287_));
 XOR2_X1 _29254_ (.A(_06711_),
    .B(_09712_),
    .Z(_00288_));
 XOR2_X2 _29255_ (.A(net794),
    .B(_10439_),
    .Z(_00241_));
 XOR2_X2 _29256_ (.A(net798),
    .B(net583),
    .Z(_00242_));
 XOR2_X2 _29257_ (.A(_06637_),
    .B(_10550_),
    .Z(_00243_));
 XOR2_X1 _29258_ (.A(_06656_),
    .B(_10535_),
    .Z(_00244_));
 XOR2_X1 _29259_ (.A(_06672_),
    .B(_10527_),
    .Z(_00245_));
 XOR2_X1 _29260_ (.A(_06687_),
    .B(_10516_),
    .Z(_00246_));
 XOR2_X1 _29261_ (.A(_06696_),
    .B(_10505_),
    .Z(_00247_));
 XOR2_X2 _29262_ (.A(_06710_),
    .B(_10432_),
    .Z(_00248_));
 XOR2_X1 _29263_ (.A(net788),
    .B(net578),
    .Z(_00209_));
 XOR2_X1 _29264_ (.A(_06619_),
    .B(net657),
    .Z(_00210_));
 XOR2_X1 _29265_ (.A(_06635_),
    .B(_11219_),
    .Z(_00211_));
 XOR2_X1 _29266_ (.A(_06654_),
    .B(_11245_),
    .Z(_00212_));
 XOR2_X1 _29267_ (.A(_06670_),
    .B(_11265_),
    .Z(_00213_));
 XOR2_X1 _29268_ (.A(_06685_),
    .B(_11202_),
    .Z(_00214_));
 XOR2_X1 _29269_ (.A(_06699_),
    .B(_11187_),
    .Z(_00215_));
 XOR2_X1 _29270_ (.A(_06708_),
    .B(_11119_),
    .Z(_00216_));
 XOR2_X2 _29271_ (.A(_06241_),
    .B(_08986_),
    .Z(_00177_));
 XOR2_X1 _29272_ (.A(_06255_),
    .B(net630),
    .Z(_00178_));
 XOR2_X2 _29273_ (.A(net1003),
    .B(_09040_),
    .Z(_00179_));
 XOR2_X1 _29274_ (.A(_06221_),
    .B(_09092_),
    .Z(_00180_));
 XOR2_X1 _29275_ (.A(_06281_),
    .B(_09161_),
    .Z(_00181_));
 XOR2_X1 _29276_ (.A(_06269_),
    .B(_09070_),
    .Z(_00182_));
 XOR2_X1 _29277_ (.A(_06575_),
    .B(_09066_),
    .Z(_00183_));
 XOR2_X1 _29278_ (.A(_06587_),
    .B(_08979_),
    .Z(_00184_));
 XOR2_X2 _29279_ (.A(_06242_),
    .B(\sa11_sr[0] ),
    .Z(_00273_));
 XOR2_X1 _29280_ (.A(_06256_),
    .B(\sa11_sr[1] ),
    .Z(_00274_));
 XOR2_X1 _29281_ (.A(_06297_),
    .B(_09762_),
    .Z(_00275_));
 XOR2_X1 _29282_ (.A(_06222_),
    .B(_09839_),
    .Z(_00276_));
 XOR2_X1 _29283_ (.A(_06282_),
    .B(_09808_),
    .Z(_00277_));
 XOR2_X2 _29284_ (.A(_06270_),
    .B(_09785_),
    .Z(_00278_));
 XOR2_X1 _29285_ (.A(_06576_),
    .B(_09786_),
    .Z(_00279_));
 XOR2_X1 _29286_ (.A(_06588_),
    .B(\sa11_sr[7] ),
    .Z(_00280_));
 XOR2_X2 _29287_ (.A(_06247_),
    .B(net529),
    .Z(_00233_));
 XOR2_X1 _29288_ (.A(_06260_),
    .B(\sa12_sr[1] ),
    .Z(_00234_));
 XOR2_X2 _29289_ (.A(_06299_),
    .B(_10478_),
    .Z(_00235_));
 XOR2_X1 _29290_ (.A(_06228_),
    .B(_10539_),
    .Z(_00236_));
 XOR2_X2 _29291_ (.A(_06284_),
    .B(_10526_),
    .Z(_00237_));
 XOR2_X1 _29292_ (.A(_06272_),
    .B(_10515_),
    .Z(_00238_));
 XOR2_X1 _29293_ (.A(_06578_),
    .B(_10502_),
    .Z(_00239_));
 XOR2_X1 _29294_ (.A(_06590_),
    .B(net551),
    .Z(_00240_));
 XOR2_X1 _29295_ (.A(net569),
    .B(\sa10_sub[0] ),
    .Z(_00201_));
 XOR2_X1 _29296_ (.A(\u0.tmp_w[17] ),
    .B(_11114_),
    .Z(_00202_));
 XOR2_X1 _29297_ (.A(_06295_),
    .B(_11158_),
    .Z(_00203_));
 XOR2_X2 _29298_ (.A(_06229_),
    .B(_11223_),
    .Z(_00204_));
 XOR2_X1 _29299_ (.A(_06285_),
    .B(_11249_),
    .Z(_00205_));
 XOR2_X2 _29300_ (.A(_06268_),
    .B(_11201_),
    .Z(_00206_));
 XOR2_X1 _29301_ (.A(_06574_),
    .B(_11186_),
    .Z(_00207_));
 XOR2_X1 _29302_ (.A(_06586_),
    .B(_11120_),
    .Z(_00208_));
 XOR2_X2 _29303_ (.A(_06450_),
    .B(net1103),
    .Z(_00169_));
 XOR2_X2 _29304_ (.A(_06465_),
    .B(net696),
    .Z(_00170_));
 XOR2_X2 _29305_ (.A(_06480_),
    .B(_09041_),
    .Z(_00171_));
 XOR2_X2 _29306_ (.A(_06510_),
    .B(_09089_),
    .Z(_00172_));
 XOR2_X2 _29307_ (.A(_06527_),
    .B(_09187_),
    .Z(_00173_));
 XOR2_X1 _29308_ (.A(_06542_),
    .B(_09165_),
    .Z(_00174_));
 XOR2_X2 _29309_ (.A(_06555_),
    .B(_09067_),
    .Z(_00175_));
 XOR2_X2 _29310_ (.A(_06564_),
    .B(_09151_),
    .Z(_00176_));
 XOR2_X1 _29311_ (.A(_06451_),
    .B(\sa21_sr[0] ),
    .Z(_00257_));
 XOR2_X2 _29312_ (.A(_06466_),
    .B(net643),
    .Z(_00258_));
 XOR2_X1 _29313_ (.A(_06483_),
    .B(_09763_),
    .Z(_00259_));
 XOR2_X1 _29314_ (.A(_06511_),
    .B(_09836_),
    .Z(_00260_));
 XOR2_X1 _29315_ (.A(_06528_),
    .B(_09869_),
    .Z(_00261_));
 XOR2_X2 _29316_ (.A(_06543_),
    .B(_09814_),
    .Z(_00262_));
 XOR2_X1 _29317_ (.A(_06556_),
    .B(_09787_),
    .Z(_00263_));
 XOR2_X2 _29318_ (.A(_06565_),
    .B(_09796_),
    .Z(_00264_));
 XOR2_X2 _29319_ (.A(_06456_),
    .B(net596),
    .Z(_00225_));
 XOR2_X1 _29320_ (.A(_06470_),
    .B(net558),
    .Z(_00226_));
 XOR2_X2 _29321_ (.A(_06482_),
    .B(_10479_),
    .Z(_00227_));
 XOR2_X1 _29322_ (.A(_06516_),
    .B(_10551_),
    .Z(_00228_));
 XOR2_X1 _29323_ (.A(_06532_),
    .B(_10536_),
    .Z(_00229_));
 XOR2_X1 _29324_ (.A(_06545_),
    .B(_10523_),
    .Z(_00230_));
 XOR2_X1 _29325_ (.A(_06558_),
    .B(_10513_),
    .Z(_00231_));
 XOR2_X1 _29326_ (.A(_06567_),
    .B(_10503_),
    .Z(_00232_));
 XOR2_X2 _29327_ (.A(_06457_),
    .B(_11136_),
    .Z(_00193_));
 XOR2_X2 _29328_ (.A(net1048),
    .B(net973),
    .Z(_00194_));
 XOR2_X2 _29329_ (.A(_06479_),
    .B(_11159_),
    .Z(_00195_));
 XOR2_X2 _29330_ (.A(_06517_),
    .B(_11220_),
    .Z(_00196_));
 XOR2_X2 _29331_ (.A(_06533_),
    .B(_11246_),
    .Z(_00197_));
 XOR2_X2 _29332_ (.A(_06546_),
    .B(_11261_),
    .Z(_00198_));
 XOR2_X1 _29333_ (.A(_06554_),
    .B(_11199_),
    .Z(_00199_));
 XOR2_X2 _29334_ (.A(_06563_),
    .B(_11183_),
    .Z(_00200_));
 XOR2_X1 _29335_ (.A(_06325_),
    .B(\sa30_sr[0] ),
    .Z(_00161_));
 XOR2_X1 _29336_ (.A(_06340_),
    .B(_08987_),
    .Z(_00162_));
 XOR2_X1 _29337_ (.A(_06355_),
    .B(_09037_),
    .Z(_00163_));
 XOR2_X1 _29338_ (.A(_06386_),
    .B(_09094_),
    .Z(_00164_));
 XOR2_X1 _29339_ (.A(_06403_),
    .B(_09190_),
    .Z(_00165_));
 XOR2_X1 _29340_ (.A(_06417_),
    .B(_09166_),
    .Z(_00166_));
 XOR2_X2 _29341_ (.A(_06431_),
    .B(_09071_),
    .Z(_00167_));
 XOR2_X1 _29342_ (.A(_06439_),
    .B(_09152_),
    .Z(_00168_));
 XOR2_X1 _29343_ (.A(_06326_),
    .B(net641),
    .Z(_00249_));
 XOR2_X1 _29344_ (.A(_06341_),
    .B(net754),
    .Z(_00250_));
 XOR2_X1 _29345_ (.A(_06356_),
    .B(_09759_),
    .Z(_00251_));
 XOR2_X1 _29346_ (.A(_06387_),
    .B(_09841_),
    .Z(_00252_));
 XOR2_X1 _29347_ (.A(_06404_),
    .B(_09872_),
    .Z(_00253_));
 XOR2_X1 _29348_ (.A(_06418_),
    .B(_09809_),
    .Z(_00254_));
 XOR2_X1 _29349_ (.A(_06432_),
    .B(_09790_),
    .Z(_00255_));
 XOR2_X1 _29350_ (.A(_06440_),
    .B(_09799_),
    .Z(_00256_));
 XOR2_X1 _29351_ (.A(_06330_),
    .B(_10453_),
    .Z(_00217_));
 XOR2_X1 _29352_ (.A(_06346_),
    .B(net544),
    .Z(_00218_));
 XOR2_X1 _29353_ (.A(_06358_),
    .B(_10475_),
    .Z(_00219_));
 XOR2_X2 _29354_ (.A(_06392_),
    .B(_10554_),
    .Z(_00220_));
 XOR2_X1 _29355_ (.A(_06406_),
    .B(_10541_),
    .Z(_00221_));
 XOR2_X1 _29356_ (.A(_06420_),
    .B(_10524_),
    .Z(_00222_));
 XOR2_X1 _29357_ (.A(_06434_),
    .B(_10512_),
    .Z(_00223_));
 XOR2_X1 _29358_ (.A(_06442_),
    .B(_10506_),
    .Z(_00224_));
 XOR2_X1 _29359_ (.A(net1020),
    .B(_11135_),
    .Z(_00265_));
 XOR2_X1 _29360_ (.A(net1018),
    .B(net971),
    .Z(_00266_));
 XOR2_X2 _29361_ (.A(_06354_),
    .B(_11164_),
    .Z(_00267_));
 XOR2_X2 _29362_ (.A(_06393_),
    .B(_11225_),
    .Z(_00268_));
 XOR2_X2 _29363_ (.A(_06407_),
    .B(_11250_),
    .Z(_00269_));
 XOR2_X1 _29364_ (.A(_06416_),
    .B(_11262_),
    .Z(_00270_));
 XOR2_X1 _29365_ (.A(_06430_),
    .B(_11198_),
    .Z(_00271_));
 XOR2_X1 _29366_ (.A(\u0.tmp_w[7] ),
    .B(_11184_),
    .Z(_00272_));
 MUX2_X1 _29367_ (.A(\text_in_r[0] ),
    .B(net228),
    .S(_06776_),
    .Z(_00489_));
 MUX2_X1 _29368_ (.A(\text_in_r[100] ),
    .B(net229),
    .S(_06776_),
    .Z(_00490_));
 MUX2_X1 _29369_ (.A(\text_in_r[101] ),
    .B(net230),
    .S(_06776_),
    .Z(_00491_));
 MUX2_X1 _29370_ (.A(\text_in_r[102] ),
    .B(net231),
    .S(_06776_),
    .Z(_00492_));
 BUF_X4 _29371_ (.A(_06771_),
    .Z(_06177_));
 MUX2_X1 _29372_ (.A(\text_in_r[103] ),
    .B(net232),
    .S(_06177_),
    .Z(_00493_));
 MUX2_X1 _29373_ (.A(\text_in_r[104] ),
    .B(net233),
    .S(_06177_),
    .Z(_00494_));
 MUX2_X1 _29374_ (.A(\text_in_r[105] ),
    .B(net234),
    .S(_06177_),
    .Z(_00495_));
 MUX2_X1 _29375_ (.A(\text_in_r[106] ),
    .B(net235),
    .S(_06177_),
    .Z(_00496_));
 MUX2_X1 _29376_ (.A(\text_in_r[107] ),
    .B(net236),
    .S(_06177_),
    .Z(_00497_));
 MUX2_X1 _29377_ (.A(\text_in_r[108] ),
    .B(net237),
    .S(_06177_),
    .Z(_00498_));
 MUX2_X1 _29378_ (.A(\text_in_r[109] ),
    .B(net238),
    .S(_06177_),
    .Z(_00499_));
 MUX2_X1 _29379_ (.A(\text_in_r[10] ),
    .B(net239),
    .S(_06177_),
    .Z(_00500_));
 MUX2_X1 _29380_ (.A(\text_in_r[110] ),
    .B(net240),
    .S(_06177_),
    .Z(_00501_));
 MUX2_X1 _29381_ (.A(\text_in_r[111] ),
    .B(net241),
    .S(_06177_),
    .Z(_00502_));
 BUF_X4 _29382_ (.A(_06771_),
    .Z(_06178_));
 MUX2_X1 _29383_ (.A(\text_in_r[112] ),
    .B(net242),
    .S(_06178_),
    .Z(_00503_));
 MUX2_X1 _29384_ (.A(\text_in_r[113] ),
    .B(net243),
    .S(_06178_),
    .Z(_00504_));
 MUX2_X1 _29385_ (.A(\text_in_r[114] ),
    .B(net244),
    .S(_06178_),
    .Z(_00505_));
 MUX2_X1 _29386_ (.A(\text_in_r[115] ),
    .B(net245),
    .S(_06178_),
    .Z(_00506_));
 MUX2_X1 _29387_ (.A(\text_in_r[116] ),
    .B(net246),
    .S(_06178_),
    .Z(_00507_));
 MUX2_X1 _29388_ (.A(\text_in_r[117] ),
    .B(net247),
    .S(_06178_),
    .Z(_00508_));
 MUX2_X1 _29389_ (.A(\text_in_r[118] ),
    .B(net248),
    .S(_06178_),
    .Z(_00509_));
 MUX2_X1 _29390_ (.A(\text_in_r[119] ),
    .B(net249),
    .S(_06178_),
    .Z(_00510_));
 MUX2_X1 _29391_ (.A(\text_in_r[11] ),
    .B(net250),
    .S(_06178_),
    .Z(_00511_));
 MUX2_X1 _29392_ (.A(\text_in_r[120] ),
    .B(net251),
    .S(_06178_),
    .Z(_00512_));
 BUF_X8 _29393_ (.A(_06401_),
    .Z(_06179_));
 BUF_X4 _29394_ (.A(_06179_),
    .Z(_06180_));
 MUX2_X1 _29395_ (.A(\text_in_r[121] ),
    .B(net252),
    .S(_06180_),
    .Z(_00513_));
 MUX2_X1 _29396_ (.A(\text_in_r[122] ),
    .B(net253),
    .S(_06180_),
    .Z(_00514_));
 MUX2_X1 _29397_ (.A(\text_in_r[123] ),
    .B(net254),
    .S(_06180_),
    .Z(_00515_));
 MUX2_X1 _29398_ (.A(\text_in_r[124] ),
    .B(net255),
    .S(_06180_),
    .Z(_00516_));
 MUX2_X1 _29399_ (.A(\text_in_r[125] ),
    .B(net256),
    .S(_06180_),
    .Z(_00517_));
 MUX2_X1 _29400_ (.A(\text_in_r[126] ),
    .B(net257),
    .S(_06180_),
    .Z(_00518_));
 MUX2_X1 _29401_ (.A(\text_in_r[127] ),
    .B(net258),
    .S(_06180_),
    .Z(_00519_));
 MUX2_X1 _29402_ (.A(\text_in_r[12] ),
    .B(net259),
    .S(_06180_),
    .Z(_00520_));
 MUX2_X1 _29403_ (.A(\text_in_r[13] ),
    .B(net260),
    .S(_06180_),
    .Z(_00521_));
 MUX2_X1 _29404_ (.A(\text_in_r[14] ),
    .B(net261),
    .S(_06180_),
    .Z(_00522_));
 BUF_X4 _29405_ (.A(_06179_),
    .Z(_06181_));
 MUX2_X1 _29406_ (.A(\text_in_r[15] ),
    .B(net262),
    .S(_06181_),
    .Z(_00523_));
 MUX2_X1 _29407_ (.A(\text_in_r[16] ),
    .B(net263),
    .S(_06181_),
    .Z(_00524_));
 MUX2_X1 _29408_ (.A(\text_in_r[17] ),
    .B(net264),
    .S(_06181_),
    .Z(_00525_));
 MUX2_X1 _29409_ (.A(\text_in_r[18] ),
    .B(net265),
    .S(_06181_),
    .Z(_00526_));
 MUX2_X1 _29410_ (.A(_13936_),
    .B(net266),
    .S(_06181_),
    .Z(_00527_));
 MUX2_X1 _29411_ (.A(\text_in_r[1] ),
    .B(net267),
    .S(_06181_),
    .Z(_00528_));
 MUX2_X1 _29412_ (.A(\text_in_r[20] ),
    .B(net268),
    .S(_06181_),
    .Z(_00529_));
 MUX2_X1 _29413_ (.A(\text_in_r[21] ),
    .B(net269),
    .S(_06181_),
    .Z(_00530_));
 MUX2_X1 _29414_ (.A(\text_in_r[22] ),
    .B(net270),
    .S(_06181_),
    .Z(_00531_));
 MUX2_X1 _29415_ (.A(\text_in_r[23] ),
    .B(net271),
    .S(_06181_),
    .Z(_00532_));
 BUF_X4 _29416_ (.A(_06179_),
    .Z(_06182_));
 MUX2_X1 _29417_ (.A(\text_in_r[24] ),
    .B(net272),
    .S(_06182_),
    .Z(_00533_));
 MUX2_X1 _29418_ (.A(\text_in_r[25] ),
    .B(net273),
    .S(_06182_),
    .Z(_00534_));
 MUX2_X1 _29419_ (.A(\text_in_r[26] ),
    .B(net274),
    .S(_06182_),
    .Z(_00535_));
 MUX2_X1 _29420_ (.A(\text_in_r[27] ),
    .B(net275),
    .S(_06182_),
    .Z(_00536_));
 MUX2_X1 _29421_ (.A(\text_in_r[28] ),
    .B(net276),
    .S(_06182_),
    .Z(_00537_));
 MUX2_X1 _29422_ (.A(\text_in_r[29] ),
    .B(net277),
    .S(_06182_),
    .Z(_00538_));
 MUX2_X1 _29423_ (.A(\text_in_r[2] ),
    .B(net278),
    .S(_06182_),
    .Z(_00539_));
 MUX2_X1 _29424_ (.A(\text_in_r[30] ),
    .B(net279),
    .S(_06182_),
    .Z(_00540_));
 MUX2_X1 _29425_ (.A(\text_in_r[31] ),
    .B(net280),
    .S(_06182_),
    .Z(_00541_));
 MUX2_X1 _29426_ (.A(\text_in_r[32] ),
    .B(net281),
    .S(_06182_),
    .Z(_00542_));
 BUF_X4 _29427_ (.A(_06179_),
    .Z(_06183_));
 MUX2_X1 _29428_ (.A(\text_in_r[33] ),
    .B(net282),
    .S(_06183_),
    .Z(_00543_));
 MUX2_X1 _29429_ (.A(\text_in_r[34] ),
    .B(net283),
    .S(_06183_),
    .Z(_00544_));
 MUX2_X1 _29430_ (.A(_04941_),
    .B(net284),
    .S(_06183_),
    .Z(_00545_));
 MUX2_X1 _29431_ (.A(\text_in_r[36] ),
    .B(net285),
    .S(_06183_),
    .Z(_00546_));
 MUX2_X1 _29432_ (.A(\text_in_r[37] ),
    .B(net286),
    .S(_06183_),
    .Z(_00547_));
 MUX2_X1 _29433_ (.A(\text_in_r[38] ),
    .B(net287),
    .S(_06183_),
    .Z(_00548_));
 MUX2_X1 _29434_ (.A(\text_in_r[39] ),
    .B(net288),
    .S(_06183_),
    .Z(_00549_));
 MUX2_X1 _29435_ (.A(\text_in_r[3] ),
    .B(net289),
    .S(_06183_),
    .Z(_00550_));
 MUX2_X1 _29436_ (.A(\text_in_r[40] ),
    .B(net290),
    .S(_06183_),
    .Z(_00551_));
 MUX2_X1 _29437_ (.A(\text_in_r[41] ),
    .B(net291),
    .S(_06183_),
    .Z(_00552_));
 BUF_X4 _29438_ (.A(_06179_),
    .Z(_06184_));
 MUX2_X1 _29439_ (.A(\text_in_r[42] ),
    .B(net292),
    .S(_06184_),
    .Z(_00553_));
 MUX2_X1 _29440_ (.A(_02333_),
    .B(net293),
    .S(_06184_),
    .Z(_00554_));
 MUX2_X1 _29441_ (.A(\text_in_r[44] ),
    .B(net294),
    .S(_06184_),
    .Z(_00555_));
 MUX2_X1 _29442_ (.A(\text_in_r[45] ),
    .B(net295),
    .S(_06184_),
    .Z(_00556_));
 MUX2_X1 _29443_ (.A(\text_in_r[46] ),
    .B(net296),
    .S(_06184_),
    .Z(_00557_));
 MUX2_X1 _29444_ (.A(\text_in_r[47] ),
    .B(net297),
    .S(_06184_),
    .Z(_00558_));
 MUX2_X1 _29445_ (.A(\text_in_r[48] ),
    .B(net298),
    .S(_06184_),
    .Z(_00559_));
 MUX2_X1 _29446_ (.A(\text_in_r[49] ),
    .B(net299),
    .S(_06184_),
    .Z(_00560_));
 MUX2_X1 _29447_ (.A(\text_in_r[4] ),
    .B(net300),
    .S(_06184_),
    .Z(_00561_));
 MUX2_X1 _29448_ (.A(\text_in_r[50] ),
    .B(net301),
    .S(_06184_),
    .Z(_00562_));
 BUF_X4 _29449_ (.A(_06179_),
    .Z(_06185_));
 MUX2_X1 _29450_ (.A(\text_in_r[51] ),
    .B(net302),
    .S(_06185_),
    .Z(_00563_));
 MUX2_X1 _29451_ (.A(\text_in_r[52] ),
    .B(net303),
    .S(_06185_),
    .Z(_00564_));
 MUX2_X1 _29452_ (.A(\text_in_r[53] ),
    .B(net304),
    .S(_06185_),
    .Z(_00565_));
 MUX2_X1 _29453_ (.A(\text_in_r[54] ),
    .B(net305),
    .S(_06185_),
    .Z(_00566_));
 MUX2_X1 _29454_ (.A(\text_in_r[55] ),
    .B(net306),
    .S(_06185_),
    .Z(_00567_));
 MUX2_X1 _29455_ (.A(\text_in_r[56] ),
    .B(net307),
    .S(_06185_),
    .Z(_00568_));
 MUX2_X1 _29456_ (.A(\text_in_r[57] ),
    .B(net308),
    .S(_06185_),
    .Z(_00569_));
 MUX2_X1 _29457_ (.A(\text_in_r[58] ),
    .B(net309),
    .S(_06185_),
    .Z(_00570_));
 MUX2_X1 _29458_ (.A(\text_in_r[59] ),
    .B(net310),
    .S(_06185_),
    .Z(_00571_));
 MUX2_X1 _29459_ (.A(\text_in_r[5] ),
    .B(net311),
    .S(_06185_),
    .Z(_00572_));
 BUF_X4 _29460_ (.A(_06179_),
    .Z(_06186_));
 MUX2_X1 _29461_ (.A(\text_in_r[60] ),
    .B(net312),
    .S(_06186_),
    .Z(_00573_));
 MUX2_X1 _29462_ (.A(\text_in_r[61] ),
    .B(net313),
    .S(_06186_),
    .Z(_00574_));
 MUX2_X1 _29463_ (.A(\text_in_r[62] ),
    .B(net314),
    .S(_06186_),
    .Z(_00575_));
 MUX2_X1 _29464_ (.A(\text_in_r[63] ),
    .B(net315),
    .S(_06186_),
    .Z(_00576_));
 MUX2_X1 _29465_ (.A(\text_in_r[64] ),
    .B(net316),
    .S(_06186_),
    .Z(_00577_));
 MUX2_X1 _29466_ (.A(\text_in_r[65] ),
    .B(net317),
    .S(_06186_),
    .Z(_00578_));
 MUX2_X1 _29467_ (.A(\text_in_r[66] ),
    .B(net318),
    .S(_06186_),
    .Z(_00579_));
 MUX2_X1 _29468_ (.A(\text_in_r[67] ),
    .B(net319),
    .S(_06186_),
    .Z(_00580_));
 MUX2_X1 _29469_ (.A(\text_in_r[68] ),
    .B(net320),
    .S(_06186_),
    .Z(_00581_));
 MUX2_X1 _29470_ (.A(\text_in_r[69] ),
    .B(net321),
    .S(_06186_),
    .Z(_00582_));
 BUF_X4 _29471_ (.A(_06179_),
    .Z(_06187_));
 MUX2_X1 _29472_ (.A(\text_in_r[6] ),
    .B(net322),
    .S(_06187_),
    .Z(_00583_));
 MUX2_X1 _29473_ (.A(\text_in_r[70] ),
    .B(net323),
    .S(_06187_),
    .Z(_00584_));
 MUX2_X1 _29474_ (.A(\text_in_r[71] ),
    .B(net324),
    .S(_06187_),
    .Z(_00585_));
 MUX2_X1 _29475_ (.A(\text_in_r[72] ),
    .B(net325),
    .S(_06187_),
    .Z(_00586_));
 MUX2_X1 _29476_ (.A(\text_in_r[73] ),
    .B(net326),
    .S(_06187_),
    .Z(_00587_));
 MUX2_X1 _29477_ (.A(\text_in_r[74] ),
    .B(net327),
    .S(_06187_),
    .Z(_00588_));
 MUX2_X1 _29478_ (.A(\text_in_r[75] ),
    .B(net328),
    .S(_06187_),
    .Z(_00589_));
 MUX2_X1 _29479_ (.A(\text_in_r[76] ),
    .B(net329),
    .S(_06187_),
    .Z(_00590_));
 MUX2_X1 _29480_ (.A(\text_in_r[77] ),
    .B(net330),
    .S(_06187_),
    .Z(_00591_));
 MUX2_X1 _29481_ (.A(\text_in_r[78] ),
    .B(net331),
    .S(_06187_),
    .Z(_00592_));
 BUF_X4 _29482_ (.A(_06179_),
    .Z(_06188_));
 MUX2_X1 _29483_ (.A(\text_in_r[79] ),
    .B(net332),
    .S(_06188_),
    .Z(_00593_));
 MUX2_X1 _29484_ (.A(\text_in_r[7] ),
    .B(net333),
    .S(_06188_),
    .Z(_00594_));
 MUX2_X1 _29485_ (.A(\text_in_r[80] ),
    .B(net334),
    .S(_06188_),
    .Z(_00595_));
 MUX2_X1 _29486_ (.A(\text_in_r[81] ),
    .B(net335),
    .S(_06188_),
    .Z(_00596_));
 MUX2_X1 _29487_ (.A(\text_in_r[82] ),
    .B(net336),
    .S(_06188_),
    .Z(_00597_));
 MUX2_X1 _29488_ (.A(\text_in_r[83] ),
    .B(net337),
    .S(_06188_),
    .Z(_00598_));
 MUX2_X1 _29489_ (.A(\text_in_r[84] ),
    .B(net338),
    .S(_06188_),
    .Z(_00599_));
 MUX2_X1 _29490_ (.A(\text_in_r[85] ),
    .B(net339),
    .S(_06188_),
    .Z(_00600_));
 MUX2_X1 _29491_ (.A(\text_in_r[86] ),
    .B(net340),
    .S(_06188_),
    .Z(_00601_));
 MUX2_X1 _29492_ (.A(\text_in_r[87] ),
    .B(net341),
    .S(_06188_),
    .Z(_00602_));
 BUF_X4 _29493_ (.A(_06179_),
    .Z(_06189_));
 MUX2_X1 _29494_ (.A(\text_in_r[88] ),
    .B(net342),
    .S(_06189_),
    .Z(_00603_));
 MUX2_X1 _29495_ (.A(\text_in_r[89] ),
    .B(net343),
    .S(_06189_),
    .Z(_00604_));
 MUX2_X1 _29496_ (.A(\text_in_r[8] ),
    .B(net344),
    .S(_06189_),
    .Z(_00605_));
 MUX2_X1 _29497_ (.A(\text_in_r[90] ),
    .B(net345),
    .S(_06189_),
    .Z(_00606_));
 MUX2_X1 _29498_ (.A(\text_in_r[91] ),
    .B(net346),
    .S(_06189_),
    .Z(_00607_));
 MUX2_X1 _29499_ (.A(\text_in_r[92] ),
    .B(net347),
    .S(_06189_),
    .Z(_00608_));
 MUX2_X1 _29500_ (.A(\text_in_r[93] ),
    .B(net348),
    .S(_06189_),
    .Z(_00609_));
 MUX2_X1 _29501_ (.A(\text_in_r[94] ),
    .B(net349),
    .S(_06189_),
    .Z(_00610_));
 MUX2_X1 _29502_ (.A(\text_in_r[95] ),
    .B(net350),
    .S(_06189_),
    .Z(_00611_));
 MUX2_X1 _29503_ (.A(\text_in_r[96] ),
    .B(net351),
    .S(_06189_),
    .Z(_00612_));
 MUX2_X1 _29504_ (.A(\text_in_r[97] ),
    .B(net352),
    .S(_06771_),
    .Z(_00613_));
 MUX2_X1 _29505_ (.A(\text_in_r[98] ),
    .B(net353),
    .S(_06771_),
    .Z(_00614_));
 MUX2_X1 _29506_ (.A(_03651_),
    .B(net354),
    .S(_06771_),
    .Z(_00615_));
 MUX2_X1 _29507_ (.A(\text_in_r[9] ),
    .B(net355),
    .S(_06771_),
    .Z(_00616_));
 INV_X1 _29508_ (.A(net227),
    .ZN(_06190_));
 INV_X1 _29509_ (.A(\dcnt[3] ),
    .ZN(_06191_));
 OR2_X1 _29510_ (.A1(\dcnt[1] ),
    .A2(_06174_),
    .ZN(_06192_));
 NOR3_X1 _29511_ (.A1(_06191_),
    .A2(_06175_),
    .A3(_06192_),
    .ZN(_06193_));
 AOI21_X1 _29512_ (.A(_06193_),
    .B1(_06192_),
    .B2(_06175_),
    .ZN(_06194_));
 NOR3_X1 _29513_ (.A1(_06772_),
    .A2(_06190_),
    .A3(_06194_),
    .ZN(_00487_));
 XNOR2_X1 _29514_ (.A(\u0.r0.rcnt[2] ),
    .B(_15330_),
    .ZN(_06195_));
 AOI21_X1 _29515_ (.A(_06776_),
    .B1(_15328_),
    .B2(_06195_),
    .ZN(_06196_));
 INV_X1 _29516_ (.A(_06196_),
    .ZN(_00617_));
 XOR2_X2 _29517_ (.A(\u0.r0.rcnt[2] ),
    .B(_15330_),
    .Z(_06197_));
 NOR2_X1 _29518_ (.A1(_06771_),
    .A2(_06197_),
    .ZN(_06198_));
 NAND3_X1 _29519_ (.A1(\u0.r0.rcnt[2] ),
    .A2(\u0.r0.rcnt[1] ),
    .A3(\u0.r0.rcnt[0] ),
    .ZN(_06199_));
 XOR2_X2 _29520_ (.A(\u0.r0.rcnt[3] ),
    .B(_06199_),
    .Z(_06200_));
 NAND2_X1 _29521_ (.A1(_15323_),
    .A2(_06200_),
    .ZN(_06201_));
 OAI21_X1 _29522_ (.A(_06201_),
    .B1(_06200_),
    .B2(\u0.r0.rcnt_next[1] ),
    .ZN(_06202_));
 AND2_X1 _29523_ (.A1(_06198_),
    .A2(_06202_),
    .ZN(_00618_));
 MUX2_X1 _29524_ (.A(_15323_),
    .B(_15326_),
    .S(_06200_),
    .Z(_06203_));
 AND2_X1 _29525_ (.A1(_06198_),
    .A2(_06203_),
    .ZN(_00619_));
 MUX2_X1 _29526_ (.A(_15328_),
    .B(_15324_),
    .S(_06200_),
    .Z(_06204_));
 AND2_X1 _29527_ (.A1(_06198_),
    .A2(_06204_),
    .ZN(_00620_));
 OR3_X1 _29528_ (.A1(\u0.r0.rcnt_next[1] ),
    .A2(_06197_),
    .A3(_06200_),
    .ZN(_06205_));
 NAND3_X1 _29529_ (.A1(_15328_),
    .A2(_06197_),
    .A3(_06200_),
    .ZN(_06206_));
 AOI21_X1 _29530_ (.A(_06772_),
    .B1(_06205_),
    .B2(_06206_),
    .ZN(_00621_));
 XNOR2_X1 _29531_ (.A(_06197_),
    .B(_06200_),
    .ZN(_06207_));
 AND3_X1 _29532_ (.A1(_06797_),
    .A2(_15323_),
    .A3(_06207_),
    .ZN(_00622_));
 NOR2_X1 _29533_ (.A1(_06401_),
    .A2(_06195_),
    .ZN(_00627_));
 AND2_X1 _29534_ (.A1(_06200_),
    .A2(_00627_),
    .ZN(_06208_));
 AND2_X1 _29535_ (.A1(_15326_),
    .A2(_06208_),
    .ZN(_00623_));
 AND2_X1 _29536_ (.A1(_15324_),
    .A2(_06208_),
    .ZN(_00624_));
 AND2_X1 _29537_ (.A1(_06797_),
    .A2(\u0.r0.rcnt_next[0] ),
    .ZN(_00625_));
 AND2_X1 _29538_ (.A1(_06797_),
    .A2(\u0.r0.rcnt_next[1] ),
    .ZN(_00626_));
 NOR2_X1 _29539_ (.A1(_06772_),
    .A2(_06200_),
    .ZN(_00628_));
 OAI21_X1 _29540_ (.A(_06721_),
    .B1(_06174_),
    .B2(_06176_),
    .ZN(_06209_));
 NAND2_X1 _29541_ (.A1(net227),
    .A2(_06209_),
    .ZN(_06210_));
 INV_X1 _29542_ (.A(_06210_),
    .ZN(_00485_));
 AOI21_X1 _29543_ (.A(_06771_),
    .B1(\dcnt[1] ),
    .B2(_06174_),
    .ZN(_06211_));
 NOR2_X1 _29544_ (.A1(\dcnt[3] ),
    .A2(_06175_),
    .ZN(_06212_));
 OAI21_X1 _29545_ (.A(_06211_),
    .B1(_06212_),
    .B2(_06192_),
    .ZN(_06213_));
 AND2_X1 _29546_ (.A1(net227),
    .A2(_06213_),
    .ZN(_00486_));
 NOR3_X1 _29547_ (.A1(\dcnt[1] ),
    .A2(_06174_),
    .A3(_06175_),
    .ZN(_06214_));
 OAI21_X1 _29548_ (.A(_06721_),
    .B1(_06191_),
    .B2(_06214_),
    .ZN(_06215_));
 AND2_X1 _29549_ (.A1(net227),
    .A2(_06215_),
    .ZN(_00488_));
 HA_X1 _29550_ (.A(_06868_),
    .B(_14659_),
    .CO(_14660_),
    .S(_14661_));
 HA_X1 _29551_ (.A(_06868_),
    .B(_14659_),
    .CO(_14662_),
    .S(_14663_));
 HA_X1 _29552_ (.A(_14664_),
    .B(_06868_),
    .CO(_14665_),
    .S(_14666_));
 HA_X1 _29553_ (.A(_14664_),
    .B(_06868_),
    .CO(_14667_),
    .S(_14668_));
 HA_X1 _29554_ (.A(_14669_),
    .B(_14659_),
    .CO(_14670_),
    .S(_14671_));
 HA_X1 _29555_ (.A(_14669_),
    .B(_14659_),
    .CO(_14672_),
    .S(_14673_));
 HA_X1 _29556_ (.A(_14669_),
    .B(_14664_),
    .CO(_14674_),
    .S(_14675_));
 HA_X1 _29557_ (.A(_14664_),
    .B(_14669_),
    .CO(_14676_),
    .S(_14677_));
 HA_X1 _29558_ (.A(net1205),
    .B(_14678_),
    .CO(_14679_),
    .S(_14680_));
 HA_X1 _29559_ (.A(net1205),
    .B(_14678_),
    .CO(_14681_),
    .S(_14682_));
 HA_X1 _29560_ (.A(net1205),
    .B(_14683_),
    .CO(_14684_),
    .S(_14685_));
 HA_X1 _29561_ (.A(_06868_),
    .B(_14683_),
    .CO(_14686_),
    .S(_14687_));
 HA_X1 _29562_ (.A(_14669_),
    .B(_14678_),
    .CO(_14688_),
    .S(_14689_));
 HA_X1 _29563_ (.A(_14669_),
    .B(_14678_),
    .CO(_14690_),
    .S(_14691_));
 HA_X1 _29564_ (.A(_14693_),
    .B(_14692_),
    .CO(_14694_),
    .S(_14695_));
 HA_X1 _29565_ (.A(_14692_),
    .B(_14693_),
    .CO(_14696_),
    .S(_14697_));
 HA_X1 _29566_ (.A(_14692_),
    .B(_14698_),
    .CO(_14699_),
    .S(_14700_));
 HA_X1 _29567_ (.A(_14698_),
    .B(_14692_),
    .CO(_14701_),
    .S(_14702_));
 HA_X1 _29568_ (.A(_14703_),
    .B(_14693_),
    .CO(_14704_),
    .S(_14705_));
 HA_X1 _29569_ (.A(_14703_),
    .B(_14693_),
    .CO(_14706_),
    .S(_14707_));
 HA_X1 _29570_ (.A(_14703_),
    .B(_14698_),
    .CO(_14708_),
    .S(_14709_));
 HA_X1 _29571_ (.A(_14703_),
    .B(_14698_),
    .CO(_14710_),
    .S(_14711_));
 HA_X1 _29572_ (.A(net15),
    .B(_14712_),
    .CO(_14713_),
    .S(_14714_));
 HA_X1 _29573_ (.A(net15),
    .B(_14712_),
    .CO(_14715_),
    .S(_14716_));
 HA_X1 _29574_ (.A(net15),
    .B(_14717_),
    .CO(_14718_),
    .S(_14719_));
 HA_X1 _29575_ (.A(_14692_),
    .B(_14717_),
    .CO(_14720_),
    .S(_14721_));
 HA_X1 _29576_ (.A(_14703_),
    .B(_14712_),
    .CO(_14722_),
    .S(_14723_));
 HA_X1 _29577_ (.A(_14703_),
    .B(_14712_),
    .CO(_14724_),
    .S(_14725_));
 HA_X1 _29578_ (.A(_07902_),
    .B(_14726_),
    .CO(_14728_),
    .S(_14729_));
 HA_X1 _29579_ (.A(_14726_),
    .B(_07902_),
    .CO(_14730_),
    .S(_14731_));
 HA_X1 _29580_ (.A(_14726_),
    .B(_14732_),
    .CO(_14733_),
    .S(_14734_));
 HA_X1 _29581_ (.A(_14732_),
    .B(_14726_),
    .CO(_14735_),
    .S(_14736_));
 HA_X1 _29582_ (.A(_07902_),
    .B(_14737_),
    .CO(_14738_),
    .S(_14739_));
 HA_X1 _29583_ (.A(_14737_),
    .B(_07902_),
    .CO(_14740_),
    .S(_14741_));
 HA_X1 _29584_ (.A(_14737_),
    .B(_14732_),
    .CO(_14742_),
    .S(_14743_));
 HA_X1 _29585_ (.A(_14737_),
    .B(_14732_),
    .CO(_14744_),
    .S(_14745_));
 HA_X1 _29586_ (.A(net29),
    .B(_14746_),
    .CO(_14747_),
    .S(_14748_));
 HA_X1 _29587_ (.A(_14726_),
    .B(_14746_),
    .CO(_14749_),
    .S(_14750_));
 HA_X1 _29588_ (.A(net29),
    .B(_14751_),
    .CO(_14752_),
    .S(_14753_));
 HA_X1 _29589_ (.A(net29),
    .B(_14751_),
    .CO(_14754_),
    .S(_14755_));
 HA_X1 _29590_ (.A(_14737_),
    .B(_14746_),
    .CO(_14756_),
    .S(_14757_));
 HA_X1 _29591_ (.A(_14737_),
    .B(_14746_),
    .CO(_14758_),
    .S(_14759_));
 HA_X1 _29592_ (.A(_14761_),
    .B(_14760_),
    .CO(_14762_),
    .S(_14763_));
 HA_X1 _29593_ (.A(_14760_),
    .B(_14761_),
    .CO(_14764_),
    .S(_14765_));
 HA_X1 _29594_ (.A(_14760_),
    .B(_14766_),
    .CO(_14767_),
    .S(_14768_));
 HA_X1 _29595_ (.A(_14760_),
    .B(_14766_),
    .CO(_14769_),
    .S(_14770_));
 HA_X1 _29596_ (.A(_14771_),
    .B(_14761_),
    .CO(_14772_),
    .S(_14773_));
 HA_X1 _29597_ (.A(_14771_),
    .B(_14761_),
    .CO(_14774_),
    .S(_14775_));
 HA_X1 _29598_ (.A(_14771_),
    .B(_14766_),
    .CO(_14776_),
    .S(_14777_));
 HA_X1 _29599_ (.A(_14771_),
    .B(_14766_),
    .CO(_14778_),
    .S(_14779_));
 HA_X1 _29600_ (.A(_14780_),
    .B(_14760_),
    .CO(_14781_),
    .S(_14782_));
 HA_X1 _29601_ (.A(_14780_),
    .B(_14760_),
    .CO(_14783_),
    .S(_14784_));
 HA_X1 _29602_ (.A(_14785_),
    .B(_14760_),
    .CO(_14786_),
    .S(_14787_));
 HA_X1 _29603_ (.A(_14785_),
    .B(_14760_),
    .CO(_14788_),
    .S(_14789_));
 HA_X1 _29604_ (.A(_14785_),
    .B(_14771_),
    .CO(_14790_),
    .S(_14791_));
 HA_X1 _29605_ (.A(_14785_),
    .B(_14771_),
    .CO(_14792_),
    .S(_14793_));
 HA_X1 _29606_ (.A(_14794_),
    .B(_14795_),
    .CO(_14796_),
    .S(_14797_));
 HA_X1 _29607_ (.A(_14794_),
    .B(_14795_),
    .CO(_14798_),
    .S(_14799_));
 HA_X1 _29608_ (.A(_14794_),
    .B(_14800_),
    .CO(_14801_),
    .S(_14802_));
 HA_X1 _29609_ (.A(_14803_),
    .B(_14795_),
    .CO(_14804_),
    .S(_14805_));
 HA_X1 _29610_ (.A(_14803_),
    .B(_14795_),
    .CO(_14806_),
    .S(_14807_));
 HA_X1 _29611_ (.A(_14803_),
    .B(_14800_),
    .CO(_14808_),
    .S(_14809_));
 HA_X1 _29612_ (.A(_14803_),
    .B(_14800_),
    .CO(_14810_),
    .S(_14811_));
 HA_X1 _29613_ (.A(_14812_),
    .B(_14795_),
    .CO(_14813_),
    .S(_14814_));
 HA_X1 _29614_ (.A(_14812_),
    .B(_14800_),
    .CO(_14815_),
    .S(_14816_));
 HA_X1 _29615_ (.A(_14812_),
    .B(_14800_),
    .CO(_14817_),
    .S(_14818_));
 HA_X1 _29616_ (.A(_14819_),
    .B(_14795_),
    .CO(_14820_),
    .S(_14821_));
 HA_X1 _29617_ (.A(_14819_),
    .B(_14795_),
    .CO(_14822_),
    .S(_14823_));
 HA_X1 _29618_ (.A(_14819_),
    .B(_14800_),
    .CO(_14824_),
    .S(_14825_));
 HA_X1 _29619_ (.A(_14826_),
    .B(_10003_),
    .CO(_14828_),
    .S(_14829_));
 HA_X1 _29620_ (.A(_14826_),
    .B(_10003_),
    .CO(_14830_),
    .S(_14831_));
 HA_X1 _29621_ (.A(_14826_),
    .B(_14832_),
    .CO(_14833_),
    .S(_14834_));
 HA_X1 _29622_ (.A(_14835_),
    .B(_10003_),
    .CO(_14836_),
    .S(_14837_));
 HA_X1 _29623_ (.A(_14835_),
    .B(_10003_),
    .CO(_14838_),
    .S(_14839_));
 HA_X1 _29624_ (.A(_14835_),
    .B(_14832_),
    .CO(_14840_),
    .S(_14841_));
 HA_X1 _29625_ (.A(_14835_),
    .B(_14832_),
    .CO(_14842_),
    .S(_14843_));
 HA_X1 _29626_ (.A(_14844_),
    .B(_10003_),
    .CO(_14845_),
    .S(_14846_));
 HA_X1 _29627_ (.A(_14844_),
    .B(_14832_),
    .CO(_14847_),
    .S(_14848_));
 HA_X1 _29628_ (.A(_14844_),
    .B(_14832_),
    .CO(_14849_),
    .S(_14850_));
 HA_X1 _29629_ (.A(_14851_),
    .B(net934),
    .CO(_14852_),
    .S(_14853_));
 HA_X1 _29630_ (.A(_14851_),
    .B(_10003_),
    .CO(_14854_),
    .S(_14855_));
 HA_X1 _29631_ (.A(_14851_),
    .B(_14832_),
    .CO(_14856_),
    .S(_14857_));
 HA_X1 _29632_ (.A(_14858_),
    .B(_14859_),
    .CO(_14860_),
    .S(_14861_));
 HA_X1 _29633_ (.A(_14858_),
    .B(_14859_),
    .CO(_14862_),
    .S(_14863_));
 HA_X1 _29634_ (.A(_14858_),
    .B(_14864_),
    .CO(_14865_),
    .S(_14866_));
 HA_X1 _29635_ (.A(_14867_),
    .B(_14859_),
    .CO(_14868_),
    .S(_14869_));
 HA_X1 _29636_ (.A(_14867_),
    .B(_14859_),
    .CO(_14870_),
    .S(_14871_));
 HA_X1 _29637_ (.A(_14867_),
    .B(_14864_),
    .CO(_14872_),
    .S(_14873_));
 HA_X1 _29638_ (.A(_14867_),
    .B(_14864_),
    .CO(_14874_),
    .S(_14875_));
 HA_X1 _29639_ (.A(_14876_),
    .B(_14859_),
    .CO(_14877_),
    .S(_14878_));
 HA_X1 _29640_ (.A(_14876_),
    .B(_14864_),
    .CO(_14879_),
    .S(_14880_));
 HA_X1 _29641_ (.A(_14876_),
    .B(_14864_),
    .CO(_14881_),
    .S(_14882_));
 HA_X1 _29642_ (.A(_14883_),
    .B(_14859_),
    .CO(_14884_),
    .S(_14885_));
 HA_X1 _29643_ (.A(_14883_),
    .B(_14859_),
    .CO(_14886_),
    .S(_14887_));
 HA_X1 _29644_ (.A(_14883_),
    .B(_14864_),
    .CO(_14888_),
    .S(_14889_));
 HA_X1 _29645_ (.A(_14890_),
    .B(_14891_),
    .CO(_14892_),
    .S(_14893_));
 HA_X1 _29646_ (.A(_14890_),
    .B(_14891_),
    .CO(_14894_),
    .S(_14895_));
 HA_X1 _29647_ (.A(_14890_),
    .B(_14896_),
    .CO(_14897_),
    .S(_14898_));
 HA_X1 _29648_ (.A(_14899_),
    .B(_14891_),
    .CO(_14900_),
    .S(_14901_));
 HA_X1 _29649_ (.A(_14899_),
    .B(_14891_),
    .CO(_14902_),
    .S(_14903_));
 HA_X1 _29650_ (.A(_14899_),
    .B(_14896_),
    .CO(_14904_),
    .S(_14905_));
 HA_X1 _29651_ (.A(_14899_),
    .B(_14896_),
    .CO(_14906_),
    .S(_14907_));
 HA_X1 _29652_ (.A(_14908_),
    .B(_14891_),
    .CO(_14909_),
    .S(_14910_));
 HA_X1 _29653_ (.A(_14908_),
    .B(_14896_),
    .CO(_14911_),
    .S(_14912_));
 HA_X1 _29654_ (.A(_14908_),
    .B(_14896_),
    .CO(_14913_),
    .S(_14914_));
 HA_X1 _29655_ (.A(_14915_),
    .B(_14891_),
    .CO(_14916_),
    .S(_14917_));
 HA_X1 _29656_ (.A(_14915_),
    .B(_14891_),
    .CO(_14918_),
    .S(_14919_));
 HA_X1 _29657_ (.A(_14915_),
    .B(_14896_),
    .CO(_14920_),
    .S(_14921_));
 HA_X1 _29658_ (.A(_14922_),
    .B(_12068_),
    .CO(_14924_),
    .S(_14925_));
 HA_X1 _29659_ (.A(_14922_),
    .B(_12068_),
    .CO(_14926_),
    .S(_14927_));
 HA_X1 _29660_ (.A(_14922_),
    .B(_14928_),
    .CO(_14929_),
    .S(_14930_));
 HA_X1 _29661_ (.A(_12068_),
    .B(_14931_),
    .CO(_14932_),
    .S(_14933_));
 HA_X1 _29662_ (.A(_12068_),
    .B(_14931_),
    .CO(_14934_),
    .S(_14935_));
 HA_X1 _29663_ (.A(_14931_),
    .B(_14928_),
    .CO(_14936_),
    .S(_14937_));
 HA_X1 _29664_ (.A(_14931_),
    .B(_14928_),
    .CO(_14938_),
    .S(_14939_));
 HA_X1 _29665_ (.A(_14940_),
    .B(net715),
    .CO(_14941_),
    .S(_14942_));
 HA_X1 _29666_ (.A(_14940_),
    .B(_14928_),
    .CO(_14943_),
    .S(_14944_));
 HA_X1 _29667_ (.A(_14940_),
    .B(_14928_),
    .CO(_14945_),
    .S(_14946_));
 HA_X1 _29668_ (.A(_14947_),
    .B(_12068_),
    .CO(_14948_),
    .S(_14949_));
 HA_X1 _29669_ (.A(_14947_),
    .B(_12068_),
    .CO(_14950_),
    .S(_14951_));
 HA_X1 _29670_ (.A(_14947_),
    .B(_14928_),
    .CO(_14952_),
    .S(_14953_));
 HA_X1 _29671_ (.A(_14955_),
    .B(_14954_),
    .CO(_14956_),
    .S(_14957_));
 HA_X1 _29672_ (.A(_14954_),
    .B(_14955_),
    .CO(_14958_),
    .S(_14959_));
 HA_X1 _29673_ (.A(_14960_),
    .B(_14954_),
    .CO(_14961_),
    .S(_14962_));
 HA_X1 _29674_ (.A(_14955_),
    .B(_14963_),
    .CO(_14964_),
    .S(_14965_));
 HA_X1 _29675_ (.A(_14963_),
    .B(_14955_),
    .CO(_14966_),
    .S(_14967_));
 HA_X1 _29676_ (.A(_14963_),
    .B(_14960_),
    .CO(_14968_),
    .S(_14969_));
 HA_X1 _29677_ (.A(_14960_),
    .B(_14963_),
    .CO(_14970_),
    .S(_14971_));
 HA_X1 _29678_ (.A(_14972_),
    .B(_14955_),
    .CO(_14973_),
    .S(_14974_));
 HA_X1 _29679_ (.A(_14972_),
    .B(_14960_),
    .CO(_14975_),
    .S(_14976_));
 HA_X1 _29680_ (.A(_14972_),
    .B(_14960_),
    .CO(_14977_),
    .S(_14978_));
 HA_X1 _29681_ (.A(_14979_),
    .B(_14955_),
    .CO(_14980_),
    .S(_14981_));
 HA_X1 _29682_ (.A(_14979_),
    .B(net200),
    .CO(_14982_),
    .S(_14983_));
 HA_X1 _29683_ (.A(_14979_),
    .B(_14960_),
    .CO(_14984_),
    .S(_14985_));
 HA_X1 _29684_ (.A(_14986_),
    .B(_14987_),
    .CO(_14988_),
    .S(_14989_));
 HA_X1 _29685_ (.A(_14986_),
    .B(_14987_),
    .CO(_14990_),
    .S(_14991_));
 HA_X1 _29686_ (.A(_14986_),
    .B(_14992_),
    .CO(_14993_),
    .S(_14994_));
 HA_X1 _29687_ (.A(_14995_),
    .B(_14987_),
    .CO(_14996_),
    .S(_14997_));
 HA_X1 _29688_ (.A(_14995_),
    .B(_14987_),
    .CO(_14998_),
    .S(_14999_));
 HA_X1 _29689_ (.A(_14995_),
    .B(_14992_),
    .CO(_15000_),
    .S(_15001_));
 HA_X1 _29690_ (.A(_14995_),
    .B(_14992_),
    .CO(_15002_),
    .S(_15003_));
 HA_X1 _29691_ (.A(_15004_),
    .B(_14987_),
    .CO(_15005_),
    .S(_15006_));
 HA_X1 _29692_ (.A(_15004_),
    .B(_14992_),
    .CO(_15007_),
    .S(_15008_));
 HA_X1 _29693_ (.A(_15004_),
    .B(_14992_),
    .CO(_15009_),
    .S(_15010_));
 HA_X1 _29694_ (.A(_15011_),
    .B(_14987_),
    .CO(_15012_),
    .S(_15013_));
 HA_X1 _29695_ (.A(_15011_),
    .B(_14987_),
    .CO(_15014_),
    .S(_15015_));
 HA_X1 _29696_ (.A(_15011_),
    .B(_14992_),
    .CO(_15016_),
    .S(_15017_));
 HA_X1 _29697_ (.A(_15018_),
    .B(_15019_),
    .CO(_15020_),
    .S(_15021_));
 HA_X1 _29698_ (.A(_15018_),
    .B(_15019_),
    .CO(_15022_),
    .S(_15023_));
 HA_X1 _29699_ (.A(_15018_),
    .B(_15024_),
    .CO(_15025_),
    .S(_15026_));
 HA_X1 _29700_ (.A(_15019_),
    .B(_15027_),
    .CO(_15028_),
    .S(_15029_));
 HA_X1 _29701_ (.A(_15027_),
    .B(_15019_),
    .CO(_15030_),
    .S(_15031_));
 HA_X1 _29702_ (.A(_15027_),
    .B(_15024_),
    .CO(_15032_),
    .S(_15033_));
 HA_X1 _29703_ (.A(_15024_),
    .B(_15027_),
    .CO(_15034_),
    .S(_15035_));
 HA_X1 _29704_ (.A(_15036_),
    .B(_15019_),
    .CO(_15037_),
    .S(_15038_));
 HA_X1 _29705_ (.A(_15036_),
    .B(_15024_),
    .CO(_15039_),
    .S(_15040_));
 HA_X1 _29706_ (.A(_15036_),
    .B(_15024_),
    .CO(_15041_),
    .S(_15042_));
 HA_X1 _29707_ (.A(_15043_),
    .B(_15019_),
    .CO(_15044_),
    .S(_15045_));
 HA_X1 _29708_ (.A(_15043_),
    .B(_15019_),
    .CO(_15046_),
    .S(_15047_));
 HA_X1 _29709_ (.A(_15043_),
    .B(_15024_),
    .CO(_15048_),
    .S(_15049_));
 HA_X1 _29710_ (.A(_15050_),
    .B(net566),
    .CO(_15052_),
    .S(_15053_));
 HA_X1 _29711_ (.A(_15050_),
    .B(net566),
    .CO(_15054_),
    .S(_15055_));
 HA_X1 _29712_ (.A(_15050_),
    .B(_00946_),
    .CO(_15057_),
    .S(_15058_));
 HA_X1 _29713_ (.A(_15050_),
    .B(_00946_),
    .CO(_15059_),
    .S(_15060_));
 HA_X1 _29714_ (.A(_15061_),
    .B(net566),
    .CO(_15062_),
    .S(_15063_));
 HA_X1 _29715_ (.A(_15061_),
    .B(net566),
    .CO(_15064_),
    .S(_15065_));
 HA_X1 _29716_ (.A(_00946_),
    .B(_15061_),
    .CO(_15066_),
    .S(_15067_));
 HA_X1 _29717_ (.A(_00946_),
    .B(_15061_),
    .CO(_15068_),
    .S(_15069_));
 HA_X1 _29718_ (.A(_15070_),
    .B(net836),
    .CO(_15071_),
    .S(_15072_));
 HA_X1 _29719_ (.A(_15070_),
    .B(net742),
    .CO(_15073_),
    .S(_15074_));
 HA_X1 _29720_ (.A(_15070_),
    .B(net1030),
    .CO(_15075_),
    .S(_15076_));
 HA_X1 _29721_ (.A(_15077_),
    .B(net836),
    .CO(_15078_),
    .S(_15079_));
 HA_X1 _29722_ (.A(_15077_),
    .B(net566),
    .CO(_15080_),
    .S(_15081_));
 HA_X1 _29723_ (.A(_15077_),
    .B(net741),
    .CO(_15082_),
    .S(_15083_));
 HA_X1 _29724_ (.A(_15077_),
    .B(net741),
    .CO(_15084_),
    .S(_15085_));
 HA_X1 _29725_ (.A(_15086_),
    .B(_15087_),
    .CO(_15088_),
    .S(_15089_));
 HA_X1 _29726_ (.A(_15086_),
    .B(_15087_),
    .CO(_15090_),
    .S(_15091_));
 HA_X1 _29727_ (.A(_15086_),
    .B(_15092_),
    .CO(_15093_),
    .S(_15094_));
 HA_X1 _29728_ (.A(_15086_),
    .B(_15092_),
    .CO(_15095_),
    .S(_15096_));
 HA_X1 _29729_ (.A(_15097_),
    .B(_15087_),
    .CO(_15098_),
    .S(_15099_));
 HA_X1 _29730_ (.A(_15097_),
    .B(_15087_),
    .CO(_15100_),
    .S(_15101_));
 HA_X1 _29731_ (.A(_15097_),
    .B(_15092_),
    .CO(_15102_),
    .S(_15103_));
 HA_X1 _29732_ (.A(_15097_),
    .B(_15092_),
    .CO(_15104_),
    .S(_15105_));
 HA_X1 _29733_ (.A(_15106_),
    .B(_15087_),
    .CO(_15107_),
    .S(_15108_));
 HA_X1 _29734_ (.A(_15106_),
    .B(_15092_),
    .CO(_15109_),
    .S(_15110_));
 HA_X1 _29735_ (.A(_15106_),
    .B(_15092_),
    .CO(_15111_),
    .S(_15112_));
 HA_X1 _29736_ (.A(_15113_),
    .B(_15087_),
    .CO(_15114_),
    .S(_15115_));
 HA_X1 _29737_ (.A(_15113_),
    .B(_15087_),
    .CO(_15116_),
    .S(_15117_));
 HA_X1 _29738_ (.A(_15113_),
    .B(_15092_),
    .CO(_15118_),
    .S(_15119_));
 HA_X1 _29739_ (.A(_15113_),
    .B(_15092_),
    .CO(_15120_),
    .S(_15121_));
 HA_X1 _29740_ (.A(_15122_),
    .B(_02314_),
    .CO(_15124_),
    .S(_15125_));
 HA_X1 _29741_ (.A(_15122_),
    .B(_02314_),
    .CO(_15126_),
    .S(_15127_));
 HA_X1 _29742_ (.A(_15122_),
    .B(_02279_),
    .CO(_15129_),
    .S(_15130_));
 HA_X1 _29743_ (.A(_15122_),
    .B(_02279_),
    .CO(_15131_),
    .S(_15132_));
 HA_X1 _29744_ (.A(_15133_),
    .B(_02314_),
    .CO(_15134_),
    .S(_15135_));
 HA_X1 _29745_ (.A(_15133_),
    .B(_02314_),
    .CO(_15136_),
    .S(_15137_));
 HA_X1 _29746_ (.A(_15133_),
    .B(_02279_),
    .CO(_15138_),
    .S(_15139_));
 HA_X1 _29747_ (.A(_15133_),
    .B(_02279_),
    .CO(_15140_),
    .S(_15141_));
 HA_X1 _29748_ (.A(_15142_),
    .B(net720),
    .CO(_15143_),
    .S(_15144_));
 HA_X1 _29749_ (.A(_15142_),
    .B(_02279_),
    .CO(_15145_),
    .S(_15146_));
 HA_X1 _29750_ (.A(_15142_),
    .B(_02279_),
    .CO(_15147_),
    .S(_15148_));
 HA_X1 _29751_ (.A(_15149_),
    .B(net145),
    .CO(_15150_),
    .S(_15151_));
 HA_X1 _29752_ (.A(_15149_),
    .B(_02314_),
    .CO(_15152_),
    .S(_15153_));
 HA_X1 _29753_ (.A(_15149_),
    .B(_02279_),
    .CO(_15154_),
    .S(_15155_));
 HA_X1 _29754_ (.A(_15149_),
    .B(_02279_),
    .CO(_15156_),
    .S(_15157_));
 HA_X1 _29755_ (.A(_15158_),
    .B(_15159_),
    .CO(_15160_),
    .S(_15161_));
 HA_X1 _29756_ (.A(_15158_),
    .B(_15159_),
    .CO(_15162_),
    .S(_15163_));
 HA_X1 _29757_ (.A(_15158_),
    .B(_15164_),
    .CO(_15165_),
    .S(_15166_));
 HA_X1 _29758_ (.A(_15158_),
    .B(_15164_),
    .CO(_15167_),
    .S(_15168_));
 HA_X1 _29759_ (.A(_15169_),
    .B(_15159_),
    .CO(_15170_),
    .S(_15171_));
 HA_X1 _29760_ (.A(_15169_),
    .B(_15159_),
    .CO(_15172_),
    .S(_15173_));
 HA_X1 _29761_ (.A(_15169_),
    .B(_15164_),
    .CO(_15174_),
    .S(_15175_));
 HA_X1 _29762_ (.A(_15169_),
    .B(_15164_),
    .CO(_15176_),
    .S(_15177_));
 HA_X1 _29763_ (.A(_15178_),
    .B(_15159_),
    .CO(_15179_),
    .S(_15180_));
 HA_X1 _29764_ (.A(_15178_),
    .B(_15164_),
    .CO(_15181_),
    .S(_15182_));
 HA_X1 _29765_ (.A(_15178_),
    .B(_15164_),
    .CO(_15183_),
    .S(_15184_));
 HA_X1 _29766_ (.A(_15185_),
    .B(_15159_),
    .CO(_15186_),
    .S(_15187_));
 HA_X1 _29767_ (.A(_15185_),
    .B(_15159_),
    .CO(_15188_),
    .S(_15189_));
 HA_X1 _29768_ (.A(_15185_),
    .B(_15164_),
    .CO(_15190_),
    .S(_15191_));
 HA_X1 _29769_ (.A(_15185_),
    .B(_15164_),
    .CO(_15192_),
    .S(_15193_));
 HA_X1 _29770_ (.A(_15194_),
    .B(_15195_),
    .CO(_15196_),
    .S(_15197_));
 HA_X1 _29771_ (.A(_15194_),
    .B(_15195_),
    .CO(_15198_),
    .S(_15199_));
 HA_X1 _29772_ (.A(_15194_),
    .B(_03588_),
    .CO(_15201_),
    .S(_15202_));
 HA_X1 _29773_ (.A(_15203_),
    .B(_15195_),
    .CO(_15204_),
    .S(_15205_));
 HA_X1 _29774_ (.A(_15195_),
    .B(_15203_),
    .CO(_15206_),
    .S(_15207_));
 HA_X1 _29775_ (.A(_15203_),
    .B(_03588_),
    .CO(_15208_),
    .S(_15209_));
 HA_X1 _29776_ (.A(_03588_),
    .B(_15203_),
    .CO(_15210_),
    .S(_15211_));
 HA_X1 _29777_ (.A(_15212_),
    .B(net154),
    .CO(_15213_),
    .S(_15214_));
 HA_X1 _29778_ (.A(_15212_),
    .B(_03588_),
    .CO(_15215_),
    .S(_15216_));
 HA_X1 _29779_ (.A(_15212_),
    .B(_03588_),
    .CO(_15217_),
    .S(_15218_));
 HA_X1 _29780_ (.A(_15219_),
    .B(_15195_),
    .CO(_15220_),
    .S(_15221_));
 HA_X1 _29781_ (.A(_15219_),
    .B(_15195_),
    .CO(_15222_),
    .S(_15223_));
 HA_X1 _29782_ (.A(_15219_),
    .B(_03588_),
    .CO(_15224_),
    .S(_15225_));
 HA_X1 _29783_ (.A(_15226_),
    .B(_04388_),
    .CO(_15228_),
    .S(_15229_));
 HA_X1 _29784_ (.A(_15226_),
    .B(_04388_),
    .CO(_15230_),
    .S(_15231_));
 HA_X1 _29785_ (.A(_15226_),
    .B(_15232_),
    .CO(_15233_),
    .S(_15234_));
 HA_X1 _29786_ (.A(_15235_),
    .B(_04388_),
    .CO(_15236_),
    .S(_15237_));
 HA_X1 _29787_ (.A(_15235_),
    .B(_04388_),
    .CO(_15238_),
    .S(_15239_));
 HA_X1 _29788_ (.A(_15235_),
    .B(_15232_),
    .CO(_15240_),
    .S(_15241_));
 HA_X1 _29789_ (.A(_15235_),
    .B(_15232_),
    .CO(_15242_),
    .S(_15243_));
 HA_X1 _29790_ (.A(_15244_),
    .B(_04388_),
    .CO(_15245_),
    .S(_15246_));
 HA_X1 _29791_ (.A(_15244_),
    .B(_15232_),
    .CO(_15247_),
    .S(_15248_));
 HA_X1 _29792_ (.A(_15244_),
    .B(_15232_),
    .CO(_15249_),
    .S(_15250_));
 HA_X1 _29793_ (.A(_15251_),
    .B(net1161),
    .CO(_15252_),
    .S(_15253_));
 HA_X1 _29794_ (.A(_15251_),
    .B(_04388_),
    .CO(_15254_),
    .S(_15255_));
 HA_X1 _29795_ (.A(_15251_),
    .B(_15232_),
    .CO(_15256_),
    .S(_15257_));
 HA_X1 _29796_ (.A(_15258_),
    .B(_15259_),
    .CO(_15260_),
    .S(_15261_));
 HA_X1 _29797_ (.A(_15258_),
    .B(_15259_),
    .CO(_15262_),
    .S(_15263_));
 HA_X1 _29798_ (.A(_15258_),
    .B(_15264_),
    .CO(_15265_),
    .S(_15266_));
 HA_X1 _29799_ (.A(_15267_),
    .B(_15259_),
    .CO(_15268_),
    .S(_15269_));
 HA_X1 _29800_ (.A(_15267_),
    .B(_15259_),
    .CO(_15270_),
    .S(_15271_));
 HA_X1 _29801_ (.A(_15267_),
    .B(_15264_),
    .CO(_15272_),
    .S(_15273_));
 HA_X1 _29802_ (.A(_15267_),
    .B(_15264_),
    .CO(_15274_),
    .S(_15275_));
 HA_X1 _29803_ (.A(_15276_),
    .B(_15259_),
    .CO(_15277_),
    .S(_15278_));
 HA_X1 _29804_ (.A(_15276_),
    .B(_15264_),
    .CO(_15279_),
    .S(_15280_));
 HA_X1 _29805_ (.A(_15276_),
    .B(_15264_),
    .CO(_15281_),
    .S(_15282_));
 HA_X1 _29806_ (.A(_15283_),
    .B(_15259_),
    .CO(_15284_),
    .S(_15285_));
 HA_X1 _29807_ (.A(_15283_),
    .B(_15259_),
    .CO(_15286_),
    .S(_15287_));
 HA_X1 _29808_ (.A(_15283_),
    .B(_15264_),
    .CO(_15288_),
    .S(_15289_));
 HA_X1 _29809_ (.A(_15290_),
    .B(_15291_),
    .CO(_15292_),
    .S(_15293_));
 HA_X1 _29810_ (.A(_15290_),
    .B(_15291_),
    .CO(_15294_),
    .S(_15295_));
 HA_X1 _29811_ (.A(_15290_),
    .B(_15296_),
    .CO(_15297_),
    .S(_15298_));
 HA_X1 _29812_ (.A(_15299_),
    .B(_15291_),
    .CO(_15300_),
    .S(_15301_));
 HA_X1 _29813_ (.A(_15299_),
    .B(_15291_),
    .CO(_15302_),
    .S(_15303_));
 HA_X1 _29814_ (.A(_15299_),
    .B(_15296_),
    .CO(_15304_),
    .S(_15305_));
 HA_X1 _29815_ (.A(_15299_),
    .B(_15296_),
    .CO(_15306_),
    .S(_15307_));
 HA_X1 _29816_ (.A(_15308_),
    .B(_15291_),
    .CO(_15309_),
    .S(_15310_));
 HA_X1 _29817_ (.A(_15308_),
    .B(_15296_),
    .CO(_15311_),
    .S(_15312_));
 HA_X1 _29818_ (.A(_15308_),
    .B(_15296_),
    .CO(_15313_),
    .S(_15314_));
 HA_X1 _29819_ (.A(_15315_),
    .B(_15291_),
    .CO(_15316_),
    .S(_15317_));
 HA_X1 _29820_ (.A(_15315_),
    .B(_15291_),
    .CO(_15318_),
    .S(_15319_));
 HA_X1 _29821_ (.A(_15315_),
    .B(_15296_),
    .CO(_15320_),
    .S(_15321_));
 HA_X1 _29822_ (.A(\u0.r0.rcnt_next[0] ),
    .B(_15322_),
    .CO(_15323_),
    .S(\u0.r0.rcnt_next[1] ));
 HA_X1 _29823_ (.A(\u0.r0.rcnt_next[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CO(_15324_),
    .S(_15325_));
 HA_X1 _29824_ (.A(\u0.r0.rcnt[0] ),
    .B(_15322_),
    .CO(_15326_),
    .S(_15327_));
 HA_X1 _29825_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CO(_15328_),
    .S(_15329_));
 HA_X1 _29826_ (.A(\u0.r0.rcnt[0] ),
    .B(\u0.r0.rcnt[1] ),
    .CO(_15330_),
    .S(_15331_));
 DFF_X1 \dcnt[0]$_SDFFE_PN0P_  (.D(_00485_),
    .CK(clknet_leaf_38_clk),
    .Q(\dcnt[0] ),
    .QN(_14264_));
 DFF_X1 \dcnt[1]$_SDFFE_PN0P_  (.D(_00486_),
    .CK(clknet_leaf_37_clk),
    .Q(\dcnt[1] ),
    .QN(_14263_));
 DFF_X1 \dcnt[2]$_SDFFE_PP0P_  (.D(_00487_),
    .CK(clknet_leaf_37_clk),
    .Q(\dcnt[2] ),
    .QN(_14262_));
 DFF_X1 \dcnt[3]$_SDFFE_PN0P_  (.D(_00488_),
    .CK(clknet_leaf_36_clk),
    .Q(\dcnt[3] ),
    .QN(_14265_));
 DFF_X1 \done$_DFF_P_  (.D(_00160_),
    .CK(clknet_leaf_37_clk),
    .Q(net356),
    .QN(_14266_));
 DFF_X1 \ld_r$_DFF_P_  (.D(net1239),
    .CK(clknet_leaf_78_clk),
    .Q(ld_r),
    .QN(_14267_));
 DFF_X2 \sa00_sr[0]$_DFF_P_  (.D(_00032_),
    .CK(clknet_leaf_76_clk),
    .Q(\sa00_sr[0] ),
    .QN(_14268_));
 DFF_X2 \sa00_sr[1]$_DFF_P_  (.D(_00033_),
    .CK(clknet_leaf_74_clk),
    .Q(\sa00_sr[1] ),
    .QN(_14269_));
 DFF_X1 \sa00_sr[2]$_DFF_P_  (.D(_00034_),
    .CK(clknet_leaf_75_clk),
    .Q(\sa00_sr[2] ),
    .QN(_14270_));
 DFF_X1 \sa00_sr[3]$_DFF_P_  (.D(_00035_),
    .CK(clknet_leaf_74_clk),
    .Q(\sa00_sr[3] ),
    .QN(_14271_));
 DFF_X1 \sa00_sr[4]$_DFF_P_  (.D(_00036_),
    .CK(clknet_leaf_72_clk),
    .Q(\sa00_sr[4] ),
    .QN(_14272_));
 DFF_X1 \sa00_sr[5]$_DFF_P_  (.D(_00037_),
    .CK(clknet_leaf_74_clk),
    .Q(\sa00_sr[5] ),
    .QN(_14273_));
 DFF_X1 \sa00_sr[6]$_DFF_P_  (.D(_00038_),
    .CK(clknet_leaf_74_clk),
    .Q(\sa00_sr[6] ),
    .QN(_14274_));
 DFF_X1 \sa00_sr[7]$_DFF_P_  (.D(_00039_),
    .CK(clknet_leaf_74_clk),
    .Q(\sa00_sr[7] ),
    .QN(_14275_));
 DFF_X1 \sa01_sr[0]$_DFF_P_  (.D(_00040_),
    .CK(clknet_leaf_42_clk),
    .Q(\sa01_sr[0] ),
    .QN(_14276_));
 DFF_X2 \sa01_sr[1]$_DFF_P_  (.D(_00041_),
    .CK(clknet_leaf_42_clk),
    .Q(\sa01_sr[1] ),
    .QN(_14277_));
 DFF_X1 \sa01_sr[2]$_DFF_P_  (.D(_00042_),
    .CK(clknet_leaf_43_clk),
    .Q(\sa01_sr[2] ),
    .QN(_14278_));
 DFF_X1 \sa01_sr[3]$_DFF_P_  (.D(_00043_),
    .CK(clknet_leaf_43_clk),
    .Q(\sa01_sr[3] ),
    .QN(_14279_));
 DFF_X1 \sa01_sr[4]$_DFF_P_  (.D(_00044_),
    .CK(clknet_leaf_44_clk),
    .Q(\sa01_sr[4] ),
    .QN(_14280_));
 DFF_X1 \sa01_sr[5]$_DFF_P_  (.D(_00045_),
    .CK(clknet_leaf_43_clk),
    .Q(\sa01_sr[5] ),
    .QN(_14281_));
 DFF_X1 \sa01_sr[6]$_DFF_P_  (.D(_00046_),
    .CK(clknet_leaf_44_clk),
    .Q(\sa01_sr[6] ),
    .QN(_14282_));
 DFF_X1 \sa01_sr[7]$_DFF_P_  (.D(_00047_),
    .CK(clknet_leaf_43_clk),
    .Q(\sa01_sr[7] ),
    .QN(_14283_));
 DFF_X1 \sa02_sr[0]$_DFF_P_  (.D(_00048_),
    .CK(clknet_leaf_64_clk),
    .Q(\sa02_sr[0] ),
    .QN(_14284_));
 DFF_X2 \sa02_sr[1]$_DFF_P_  (.D(_00049_),
    .CK(clknet_leaf_63_clk),
    .Q(\sa02_sr[1] ),
    .QN(_14285_));
 DFF_X1 \sa02_sr[2]$_DFF_P_  (.D(_00050_),
    .CK(clknet_leaf_45_clk),
    .Q(\sa02_sr[2] ),
    .QN(_14286_));
 DFF_X1 \sa02_sr[3]$_DFF_P_  (.D(_00051_),
    .CK(clknet_leaf_67_clk),
    .Q(\sa02_sr[3] ),
    .QN(_14287_));
 DFF_X1 \sa02_sr[4]$_DFF_P_  (.D(_00052_),
    .CK(clknet_leaf_65_clk),
    .Q(\sa02_sr[4] ),
    .QN(_14288_));
 DFF_X1 \sa02_sr[5]$_DFF_P_  (.D(_00053_),
    .CK(clknet_leaf_66_clk),
    .Q(\sa02_sr[5] ),
    .QN(_14289_));
 DFF_X1 \sa02_sr[6]$_DFF_P_  (.D(_00054_),
    .CK(clknet_leaf_64_clk),
    .Q(\sa02_sr[6] ),
    .QN(_14290_));
 DFF_X1 \sa02_sr[7]$_DFF_P_  (.D(_00055_),
    .CK(clknet_leaf_64_clk),
    .Q(\sa02_sr[7] ),
    .QN(_14291_));
 DFF_X2 \sa03_sr[0]$_DFF_P_  (.D(_00056_),
    .CK(clknet_leaf_16_clk),
    .Q(\sa03_sr[0] ),
    .QN(_14292_));
 DFF_X1 \sa03_sr[1]$_DFF_P_  (.D(_00057_),
    .CK(clknet_leaf_17_clk),
    .Q(\sa03_sr[1] ),
    .QN(_14293_));
 DFF_X1 \sa03_sr[2]$_DFF_P_  (.D(_00058_),
    .CK(clknet_leaf_17_clk),
    .Q(\sa03_sr[2] ),
    .QN(_14294_));
 DFF_X1 \sa03_sr[3]$_DFF_P_  (.D(_00059_),
    .CK(clknet_leaf_16_clk),
    .Q(\sa03_sr[3] ),
    .QN(_14295_));
 DFF_X1 \sa03_sr[4]$_DFF_P_  (.D(_00060_),
    .CK(clknet_leaf_16_clk),
    .Q(\sa03_sr[4] ),
    .QN(_14296_));
 DFF_X1 \sa03_sr[5]$_DFF_P_  (.D(_00061_),
    .CK(clknet_leaf_17_clk),
    .Q(\sa03_sr[5] ),
    .QN(_14297_));
 DFF_X1 \sa03_sr[6]$_DFF_P_  (.D(_00062_),
    .CK(clknet_leaf_16_clk),
    .Q(\sa03_sr[6] ),
    .QN(_14298_));
 DFF_X1 \sa03_sr[7]$_DFF_P_  (.D(_00063_),
    .CK(clknet_leaf_17_clk),
    .Q(\sa03_sr[7] ),
    .QN(_14299_));
 DFF_X1 \sa10_sr[0]$_DFF_P_  (.D(_00072_),
    .CK(clknet_leaf_76_clk),
    .Q(\sa10_sr[0] ),
    .QN(_14300_));
 DFF_X2 \sa10_sr[1]$_DFF_P_  (.D(_00073_),
    .CK(clknet_leaf_77_clk),
    .Q(\sa10_sr[1] ),
    .QN(_14301_));
 DFF_X1 \sa10_sr[2]$_DFF_P_  (.D(_00074_),
    .CK(clknet_leaf_77_clk),
    .Q(\sa10_sr[2] ),
    .QN(_14302_));
 DFF_X1 \sa10_sr[3]$_DFF_P_  (.D(_00075_),
    .CK(clknet_leaf_77_clk),
    .Q(\sa10_sr[3] ),
    .QN(_14303_));
 DFF_X1 \sa10_sr[4]$_DFF_P_  (.D(_00076_),
    .CK(clknet_leaf_75_clk),
    .Q(\sa10_sr[4] ),
    .QN(_14304_));
 DFF_X1 \sa10_sr[5]$_DFF_P_  (.D(_00077_),
    .CK(clknet_leaf_76_clk),
    .Q(\sa10_sr[5] ),
    .QN(_14305_));
 DFF_X1 \sa10_sr[6]$_DFF_P_  (.D(_00078_),
    .CK(clknet_leaf_75_clk),
    .Q(\sa10_sr[6] ),
    .QN(_14306_));
 DFF_X1 \sa10_sr[7]$_DFF_P_  (.D(_00079_),
    .CK(clknet_leaf_75_clk),
    .Q(\sa10_sr[7] ),
    .QN(_14307_));
 DFF_X2 \sa11_sr[0]$_DFF_P_  (.D(_00080_),
    .CK(clknet_leaf_68_clk),
    .Q(\sa11_sr[0] ),
    .QN(_14308_));
 DFF_X2 \sa11_sr[1]$_DFF_P_  (.D(net9),
    .CK(clknet_leaf_54_clk),
    .Q(\sa11_sr[1] ),
    .QN(_14309_));
 DFF_X1 \sa11_sr[2]$_DFF_P_  (.D(_00082_),
    .CK(clknet_leaf_66_clk),
    .Q(\sa11_sr[2] ),
    .QN(_14310_));
 DFF_X1 \sa11_sr[3]$_DFF_P_  (.D(_00083_),
    .CK(clknet_leaf_69_clk),
    .Q(\sa11_sr[3] ),
    .QN(_14311_));
 DFF_X1 \sa11_sr[4]$_DFF_P_  (.D(_00084_),
    .CK(clknet_leaf_66_clk),
    .Q(\sa11_sr[4] ),
    .QN(_14312_));
 DFF_X1 \sa11_sr[5]$_DFF_P_  (.D(_00085_),
    .CK(clknet_leaf_66_clk),
    .Q(\sa11_sr[5] ),
    .QN(_14313_));
 DFF_X1 \sa11_sr[6]$_DFF_P_  (.D(_00086_),
    .CK(clknet_leaf_66_clk),
    .Q(\sa11_sr[6] ),
    .QN(_14314_));
 DFF_X2 \sa11_sr[7]$_DFF_P_  (.D(_00087_),
    .CK(clknet_leaf_66_clk),
    .Q(\sa11_sr[7] ),
    .QN(_14315_));
 DFF_X2 \sa12_sr[0]$_DFF_P_  (.D(_00088_),
    .CK(clknet_leaf_79_clk),
    .Q(\sa12_sr[0] ),
    .QN(_14316_));
 DFF_X2 \sa12_sr[1]$_DFF_P_  (.D(_00089_),
    .CK(clknet_leaf_86_clk),
    .Q(\sa12_sr[1] ),
    .QN(_14317_));
 DFF_X2 \sa12_sr[2]$_DFF_P_  (.D(_00090_),
    .CK(clknet_leaf_88_clk),
    .Q(\sa12_sr[2] ),
    .QN(_14318_));
 DFF_X2 \sa12_sr[3]$_DFF_P_  (.D(_00091_),
    .CK(clknet_leaf_85_clk),
    .Q(\sa12_sr[3] ),
    .QN(_14319_));
 DFF_X1 \sa12_sr[4]$_DFF_P_  (.D(_00092_),
    .CK(clknet_leaf_3_clk),
    .Q(\sa12_sr[4] ),
    .QN(_14320_));
 DFF_X1 \sa12_sr[5]$_DFF_P_  (.D(_00093_),
    .CK(clknet_leaf_81_clk),
    .Q(\sa12_sr[5] ),
    .QN(_14321_));
 DFF_X1 \sa12_sr[6]$_DFF_P_  (.D(_00094_),
    .CK(clknet_leaf_87_clk),
    .Q(\sa12_sr[6] ),
    .QN(_14322_));
 DFF_X2 \sa12_sr[7]$_DFF_P_  (.D(_00095_),
    .CK(clknet_leaf_79_clk),
    .Q(\sa12_sr[7] ),
    .QN(_14323_));
 DFF_X2 \sa13_sr[0]$_DFF_P_  (.D(_00064_),
    .CK(clknet_leaf_1_clk),
    .Q(\sa10_sub[0] ),
    .QN(_14324_));
 DFF_X1 \sa13_sr[1]$_DFF_P_  (.D(_00065_),
    .CK(clknet_leaf_95_clk),
    .Q(\sa10_sub[1] ),
    .QN(_14325_));
 DFF_X1 \sa13_sr[2]$_DFF_P_  (.D(_00066_),
    .CK(clknet_leaf_96_clk),
    .Q(\sa10_sub[2] ),
    .QN(_14326_));
 DFF_X1 \sa13_sr[3]$_DFF_P_  (.D(_00067_),
    .CK(clknet_leaf_96_clk),
    .Q(\sa10_sub[3] ),
    .QN(_14327_));
 DFF_X1 \sa13_sr[4]$_DFF_P_  (.D(_00068_),
    .CK(clknet_leaf_96_clk),
    .Q(\sa10_sub[4] ),
    .QN(_14328_));
 DFF_X1 \sa13_sr[5]$_DFF_P_  (.D(_00069_),
    .CK(clknet_leaf_96_clk),
    .Q(\sa10_sub[5] ),
    .QN(_14329_));
 DFF_X1 \sa13_sr[6]$_DFF_P_  (.D(_00070_),
    .CK(clknet_leaf_96_clk),
    .Q(\sa10_sub[6] ),
    .QN(_14330_));
 DFF_X1 \sa13_sr[7]$_DFF_P_  (.D(_00071_),
    .CK(clknet_leaf_95_clk),
    .Q(\sa10_sub[7] ),
    .QN(_14331_));
 DFF_X1 \sa20_sr[0]$_DFF_P_  (.D(_00112_),
    .CK(clknet_leaf_74_clk),
    .Q(\sa20_sr[0] ),
    .QN(_14332_));
 DFF_X2 \sa20_sr[1]$_DFF_P_  (.D(_00113_),
    .CK(clknet_leaf_82_clk),
    .Q(\sa20_sr[1] ),
    .QN(_14333_));
 DFF_X1 \sa20_sr[2]$_DFF_P_  (.D(_00114_),
    .CK(clknet_leaf_70_clk),
    .Q(\sa20_sr[2] ),
    .QN(_14334_));
 DFF_X1 \sa20_sr[3]$_DFF_P_  (.D(_00115_),
    .CK(clknet_leaf_71_clk),
    .Q(\sa20_sr[3] ),
    .QN(_14335_));
 DFF_X1 \sa20_sr[4]$_DFF_P_  (.D(_00116_),
    .CK(clknet_leaf_71_clk),
    .Q(\sa20_sr[4] ),
    .QN(_14336_));
 DFF_X1 \sa20_sr[5]$_DFF_P_  (.D(_00117_),
    .CK(clknet_leaf_71_clk),
    .Q(\sa20_sr[5] ),
    .QN(_14337_));
 DFF_X1 \sa20_sr[6]$_DFF_P_  (.D(_00118_),
    .CK(clknet_leaf_71_clk),
    .Q(\sa20_sr[6] ),
    .QN(_14338_));
 DFF_X1 \sa20_sr[7]$_DFF_P_  (.D(_00119_),
    .CK(clknet_leaf_75_clk),
    .Q(\sa20_sr[7] ),
    .QN(_14339_));
 DFF_X2 \sa21_sr[0]$_DFF_P_  (.D(_00120_),
    .CK(clknet_leaf_11_clk),
    .Q(\sa21_sr[0] ),
    .QN(_14340_));
 DFF_X2 \sa21_sr[1]$_DFF_P_  (.D(_00121_),
    .CK(clknet_leaf_9_clk),
    .Q(\sa21_sr[1] ),
    .QN(_14341_));
 DFF_X1 \sa21_sr[2]$_DFF_P_  (.D(_00122_),
    .CK(clknet_leaf_18_clk),
    .Q(\sa21_sr[2] ),
    .QN(_14342_));
 DFF_X1 \sa21_sr[3]$_DFF_P_  (.D(_00123_),
    .CK(clknet_leaf_18_clk),
    .Q(\sa21_sr[3] ),
    .QN(_14343_));
 DFF_X1 \sa21_sr[4]$_DFF_P_  (.D(_00124_),
    .CK(clknet_leaf_1_clk),
    .Q(\sa21_sr[4] ),
    .QN(_14344_));
 DFF_X1 \sa21_sr[5]$_DFF_P_  (.D(_00125_),
    .CK(clknet_leaf_18_clk),
    .Q(\sa21_sr[5] ),
    .QN(_14345_));
 DFF_X1 \sa21_sr[6]$_DFF_P_  (.D(_00126_),
    .CK(clknet_leaf_1_clk),
    .Q(\sa21_sr[6] ),
    .QN(_14346_));
 DFF_X1 \sa21_sr[7]$_DFF_P_  (.D(_00127_),
    .CK(clknet_leaf_9_clk),
    .Q(\sa21_sr[7] ),
    .QN(_14347_));
 DFF_X2 \sa22_sr[0]$_DFF_P_  (.D(_00096_),
    .CK(clknet_leaf_58_clk),
    .Q(\sa20_sub[0] ),
    .QN(_14348_));
 DFF_X2 \sa22_sr[1]$_DFF_P_  (.D(_00097_),
    .CK(clknet_leaf_59_clk),
    .Q(\sa20_sub[1] ),
    .QN(_14349_));
 DFF_X1 \sa22_sr[2]$_DFF_P_  (.D(_00098_),
    .CK(clknet_leaf_59_clk),
    .Q(\sa20_sub[2] ),
    .QN(_14350_));
 DFF_X1 \sa22_sr[3]$_DFF_P_  (.D(_00099_),
    .CK(clknet_leaf_69_clk),
    .Q(\sa20_sub[3] ),
    .QN(_14351_));
 DFF_X1 \sa22_sr[4]$_DFF_P_  (.D(_00100_),
    .CK(clknet_leaf_59_clk),
    .Q(\sa20_sub[4] ),
    .QN(_14352_));
 DFF_X1 \sa22_sr[5]$_DFF_P_  (.D(_00101_),
    .CK(clknet_leaf_69_clk),
    .Q(\sa20_sub[5] ),
    .QN(_14353_));
 DFF_X1 \sa22_sr[6]$_DFF_P_  (.D(_00102_),
    .CK(clknet_leaf_70_clk),
    .Q(\sa20_sub[6] ),
    .QN(_14354_));
 DFF_X1 \sa22_sr[7]$_DFF_P_  (.D(_00103_),
    .CK(clknet_leaf_69_clk),
    .Q(\sa20_sub[7] ),
    .QN(_14355_));
 DFF_X1 \sa23_sr[0]$_DFF_P_  (.D(_00104_),
    .CK(clknet_leaf_11_clk),
    .Q(\sa21_sub[0] ),
    .QN(_14356_));
 DFF_X1 \sa23_sr[1]$_DFF_P_  (.D(_00105_),
    .CK(clknet_leaf_10_clk),
    .Q(\sa21_sub[1] ),
    .QN(_14357_));
 DFF_X1 \sa23_sr[2]$_DFF_P_  (.D(_00106_),
    .CK(clknet_leaf_10_clk),
    .Q(\sa21_sub[2] ),
    .QN(_14358_));
 DFF_X1 \sa23_sr[3]$_DFF_P_  (.D(_00107_),
    .CK(clknet_leaf_29_clk),
    .Q(\sa21_sub[3] ),
    .QN(_14359_));
 DFF_X1 \sa23_sr[4]$_DFF_P_  (.D(_00108_),
    .CK(clknet_leaf_10_clk),
    .Q(\sa21_sub[4] ),
    .QN(_14360_));
 DFF_X1 \sa23_sr[5]$_DFF_P_  (.D(_00109_),
    .CK(clknet_leaf_9_clk),
    .Q(\sa21_sub[5] ),
    .QN(_14361_));
 DFF_X1 \sa23_sr[6]$_DFF_P_  (.D(_00110_),
    .CK(clknet_leaf_9_clk),
    .Q(\sa21_sub[6] ),
    .QN(_14362_));
 DFF_X1 \sa23_sr[7]$_DFF_P_  (.D(_00111_),
    .CK(clknet_leaf_9_clk),
    .Q(\sa21_sub[7] ),
    .QN(_14363_));
 DFF_X2 \sa30_sr[0]$_DFF_P_  (.D(_00152_),
    .CK(clknet_leaf_23_clk),
    .Q(\sa30_sr[0] ),
    .QN(_14364_));
 DFF_X1 \sa30_sr[1]$_DFF_P_  (.D(_00153_),
    .CK(clknet_leaf_25_clk),
    .Q(\sa30_sr[1] ),
    .QN(_14365_));
 DFF_X1 \sa30_sr[2]$_DFF_P_  (.D(_00154_),
    .CK(clknet_leaf_26_clk),
    .Q(\sa30_sr[2] ),
    .QN(_14366_));
 DFF_X1 \sa30_sr[3]$_DFF_P_  (.D(_00155_),
    .CK(clknet_leaf_26_clk),
    .Q(\sa30_sr[3] ),
    .QN(_14367_));
 DFF_X1 \sa30_sr[4]$_DFF_P_  (.D(_00156_),
    .CK(clknet_leaf_26_clk),
    .Q(\sa30_sr[4] ),
    .QN(_14368_));
 DFF_X1 \sa30_sr[5]$_DFF_P_  (.D(_00157_),
    .CK(clknet_leaf_21_clk),
    .Q(\sa30_sr[5] ),
    .QN(_14369_));
 DFF_X1 \sa30_sr[6]$_DFF_P_  (.D(_00158_),
    .CK(clknet_leaf_26_clk),
    .Q(\sa30_sr[6] ),
    .QN(_14370_));
 DFF_X1 \sa30_sr[7]$_DFF_P_  (.D(_00159_),
    .CK(clknet_leaf_38_clk),
    .Q(\sa30_sr[7] ),
    .QN(_14371_));
 DFF_X2 \sa31_sr[0]$_DFF_P_  (.D(_00128_),
    .CK(clknet_leaf_52_clk),
    .Q(\sa30_sub[0] ),
    .QN(_14372_));
 DFF_X2 \sa31_sr[1]$_DFF_P_  (.D(_00129_),
    .CK(clknet_leaf_34_clk),
    .Q(\sa30_sub[1] ),
    .QN(_14373_));
 DFF_X1 \sa31_sr[2]$_DFF_P_  (.D(_00130_),
    .CK(clknet_leaf_39_clk),
    .Q(\sa30_sub[2] ),
    .QN(_14374_));
 DFF_X1 \sa31_sr[3]$_DFF_P_  (.D(_00131_),
    .CK(clknet_leaf_39_clk),
    .Q(\sa30_sub[3] ),
    .QN(_14375_));
 DFF_X1 \sa31_sr[4]$_DFF_P_  (.D(_00132_),
    .CK(clknet_leaf_34_clk),
    .Q(\sa30_sub[4] ),
    .QN(_14376_));
 DFF_X1 \sa31_sr[5]$_DFF_P_  (.D(_00133_),
    .CK(clknet_leaf_40_clk),
    .Q(\sa30_sub[5] ),
    .QN(_14377_));
 DFF_X1 \sa31_sr[6]$_DFF_P_  (.D(_00134_),
    .CK(clknet_leaf_40_clk),
    .Q(\sa30_sub[6] ),
    .QN(_14378_));
 DFF_X1 \sa31_sr[7]$_DFF_P_  (.D(_00135_),
    .CK(clknet_leaf_39_clk),
    .Q(\sa30_sub[7] ),
    .QN(_14379_));
 DFF_X1 \sa32_sr[0]$_DFF_P_  (.D(_00136_),
    .CK(clknet_leaf_44_clk),
    .Q(\sa31_sub[0] ),
    .QN(_14380_));
 DFF_X2 \sa32_sr[1]$_DFF_P_  (.D(_00137_),
    .CK(clknet_leaf_48_clk),
    .Q(\sa31_sub[1] ),
    .QN(_14381_));
 DFF_X1 \sa32_sr[2]$_DFF_P_  (.D(_00138_),
    .CK(clknet_leaf_40_clk),
    .Q(\sa31_sub[2] ),
    .QN(_14382_));
 DFF_X1 \sa32_sr[3]$_DFF_P_  (.D(_00139_),
    .CK(clknet_leaf_41_clk),
    .Q(\sa31_sub[3] ),
    .QN(_14383_));
 DFF_X1 \sa32_sr[4]$_DFF_P_  (.D(_00140_),
    .CK(clknet_leaf_41_clk),
    .Q(\sa31_sub[4] ),
    .QN(_14384_));
 DFF_X1 \sa32_sr[5]$_DFF_P_  (.D(_00141_),
    .CK(clknet_leaf_41_clk),
    .Q(\sa31_sub[5] ),
    .QN(_14385_));
 DFF_X1 \sa32_sr[6]$_DFF_P_  (.D(_00142_),
    .CK(clknet_leaf_42_clk),
    .Q(\sa31_sub[6] ),
    .QN(_14386_));
 DFF_X1 \sa32_sr[7]$_DFF_P_  (.D(_00143_),
    .CK(clknet_leaf_41_clk),
    .Q(\sa31_sub[7] ),
    .QN(_14387_));
 DFF_X1 \sa33_sr[0]$_DFF_P_  (.D(_00144_),
    .CK(clknet_leaf_29_clk),
    .Q(\sa32_sub[0] ),
    .QN(_14388_));
 DFF_X2 \sa33_sr[1]$_DFF_P_  (.D(_00145_),
    .CK(clknet_leaf_14_clk),
    .Q(\sa32_sub[1] ),
    .QN(_14389_));
 DFF_X2 \sa33_sr[2]$_DFF_P_  (.D(_00146_),
    .CK(clknet_leaf_33_clk),
    .Q(\sa32_sub[2] ),
    .QN(_14390_));
 DFF_X2 \sa33_sr[3]$_DFF_P_  (.D(_00147_),
    .CK(clknet_leaf_51_clk),
    .Q(\sa32_sub[3] ),
    .QN(_14391_));
 DFF_X1 \sa33_sr[4]$_DFF_P_  (.D(_00148_),
    .CK(clknet_leaf_35_clk),
    .Q(\sa32_sub[4] ),
    .QN(_14392_));
 DFF_X1 \sa33_sr[5]$_DFF_P_  (.D(_00149_),
    .CK(clknet_leaf_33_clk),
    .Q(\sa32_sub[5] ),
    .QN(_14393_));
 DFF_X1 \sa33_sr[6]$_DFF_P_  (.D(_00150_),
    .CK(clknet_leaf_34_clk),
    .Q(\sa32_sub[6] ),
    .QN(_14394_));
 DFF_X1 \sa33_sr[7]$_DFF_P_  (.D(_00151_),
    .CK(clknet_leaf_15_clk),
    .Q(\sa32_sub[7] ),
    .QN(_14261_));
 DFF_X1 \text_in_r[0]$_DFFE_PP_  (.D(_00489_),
    .CK(clknet_leaf_10_clk),
    .Q(\text_in_r[0] ),
    .QN(_00406_));
 DFF_X1 \text_in_r[100]$_DFFE_PP_  (.D(_00490_),
    .CK(clknet_leaf_55_clk),
    .Q(\text_in_r[100] ),
    .QN(_14260_));
 DFF_X1 \text_in_r[101]$_DFFE_PP_  (.D(_00491_),
    .CK(clknet_leaf_51_clk),
    .Q(\text_in_r[101] ),
    .QN(_14259_));
 DFF_X1 \text_in_r[102]$_DFFE_PP_  (.D(_00492_),
    .CK(clknet_leaf_56_clk),
    .Q(\text_in_r[102] ),
    .QN(_14258_));
 DFF_X1 \text_in_r[103]$_DFFE_PP_  (.D(_00493_),
    .CK(clknet_leaf_56_clk),
    .Q(\text_in_r[103] ),
    .QN(_14257_));
 DFF_X2 \text_in_r[104]$_DFFE_PP_  (.D(_00494_),
    .CK(clknet_leaf_73_clk),
    .Q(\text_in_r[104] ),
    .QN(_00465_));
 DFF_X1 \text_in_r[105]$_DFFE_PP_  (.D(_00495_),
    .CK(clknet_leaf_72_clk),
    .Q(\text_in_r[105] ),
    .QN(_00464_));
 DFF_X1 \text_in_r[106]$_DFFE_PP_  (.D(_00496_),
    .CK(clknet_leaf_29_clk),
    .Q(\text_in_r[106] ),
    .QN(_00466_));
 DFF_X2 \text_in_r[107]$_DFFE_PP_  (.D(_00497_),
    .CK(clknet_leaf_72_clk),
    .Q(\text_in_r[107] ),
    .QN(_14256_));
 DFF_X2 \text_in_r[108]$_DFFE_PP_  (.D(_00498_),
    .CK(clknet_leaf_72_clk),
    .Q(\text_in_r[108] ),
    .QN(_14255_));
 DFF_X2 \text_in_r[109]$_DFFE_PP_  (.D(_00499_),
    .CK(clknet_leaf_92_clk),
    .Q(\text_in_r[109] ),
    .QN(_14254_));
 DFF_X1 \text_in_r[10]$_DFFE_PP_  (.D(_00500_),
    .CK(clknet_leaf_5_clk),
    .Q(\text_in_r[10] ),
    .QN(_00475_));
 DFF_X1 \text_in_r[110]$_DFFE_PP_  (.D(_00501_),
    .CK(clknet_leaf_94_clk),
    .Q(\text_in_r[110] ),
    .QN(_14253_));
 DFF_X1 \text_in_r[111]$_DFFE_PP_  (.D(_00502_),
    .CK(clknet_leaf_73_clk),
    .Q(\text_in_r[111] ),
    .QN(_14252_));
 DFF_X1 \text_in_r[112]$_DFFE_PP_  (.D(_00503_),
    .CK(clknet_leaf_92_clk),
    .Q(\text_in_r[112] ),
    .QN(_00453_));
 DFF_X2 \text_in_r[113]$_DFFE_PP_  (.D(_00504_),
    .CK(clknet_leaf_92_clk),
    .Q(\text_in_r[113] ),
    .QN(_00452_));
 DFF_X2 \text_in_r[114]$_DFFE_PP_  (.D(_00505_),
    .CK(clknet_leaf_92_clk),
    .Q(\text_in_r[114] ),
    .QN(_00454_));
 DFF_X2 \text_in_r[115]$_DFFE_PP_  (.D(_00506_),
    .CK(clknet_leaf_95_clk),
    .Q(\text_in_r[115] ),
    .QN(_14251_));
 DFF_X1 \text_in_r[116]$_DFFE_PP_  (.D(_00507_),
    .CK(clknet_leaf_91_clk),
    .Q(\text_in_r[116] ),
    .QN(_14250_));
 DFF_X1 \text_in_r[117]$_DFFE_PP_  (.D(_00508_),
    .CK(clknet_leaf_84_clk),
    .Q(\text_in_r[117] ),
    .QN(_14249_));
 DFF_X1 \text_in_r[118]$_DFFE_PP_  (.D(_00509_),
    .CK(clknet_leaf_90_clk),
    .Q(\text_in_r[118] ),
    .QN(_14248_));
 DFF_X1 \text_in_r[119]$_DFFE_PP_  (.D(_00510_),
    .CK(clknet_leaf_93_clk),
    .Q(\text_in_r[119] ),
    .QN(_14247_));
 DFF_X1 \text_in_r[11]$_DFFE_PP_  (.D(_00511_),
    .CK(clknet_leaf_4_clk),
    .Q(\text_in_r[11] ),
    .QN(_14246_));
 DFF_X1 \text_in_r[120]$_DFFE_PP_  (.D(_00512_),
    .CK(clknet_leaf_91_clk),
    .Q(\text_in_r[120] ),
    .QN(_00441_));
 DFF_X1 \text_in_r[121]$_DFFE_PP_  (.D(_00513_),
    .CK(clknet_leaf_91_clk),
    .Q(\text_in_r[121] ),
    .QN(_00440_));
 DFF_X2 \text_in_r[122]$_DFFE_PP_  (.D(_00514_),
    .CK(clknet_leaf_93_clk),
    .Q(\text_in_r[122] ),
    .QN(_00442_));
 DFF_X2 \text_in_r[123]$_DFFE_PP_  (.D(_00515_),
    .CK(clknet_leaf_93_clk),
    .Q(\text_in_r[123] ),
    .QN(_14245_));
 DFF_X2 \text_in_r[124]$_DFFE_PP_  (.D(_00516_),
    .CK(clknet_leaf_73_clk),
    .Q(\text_in_r[124] ),
    .QN(_14244_));
 DFF_X2 \text_in_r[125]$_DFFE_PP_  (.D(_00517_),
    .CK(clknet_leaf_93_clk),
    .Q(\text_in_r[125] ),
    .QN(_14243_));
 DFF_X1 \text_in_r[126]$_DFFE_PP_  (.D(_00518_),
    .CK(clknet_leaf_72_clk),
    .Q(\text_in_r[126] ),
    .QN(_14242_));
 DFF_X1 \text_in_r[127]$_DFFE_PP_  (.D(_00519_),
    .CK(clknet_leaf_73_clk),
    .Q(\text_in_r[127] ),
    .QN(_14241_));
 DFF_X1 \text_in_r[12]$_DFFE_PP_  (.D(_00520_),
    .CK(clknet_leaf_4_clk),
    .Q(\text_in_r[12] ),
    .QN(_14240_));
 DFF_X1 \text_in_r[13]$_DFFE_PP_  (.D(_00521_),
    .CK(clknet_leaf_4_clk),
    .Q(\text_in_r[13] ),
    .QN(_14239_));
 DFF_X1 \text_in_r[14]$_DFFE_PP_  (.D(_00522_),
    .CK(clknet_leaf_19_clk),
    .Q(\text_in_r[14] ),
    .QN(_14238_));
 DFF_X1 \text_in_r[15]$_DFFE_PP_  (.D(_00523_),
    .CK(clknet_leaf_19_clk),
    .Q(\text_in_r[15] ),
    .QN(_14237_));
 DFF_X2 \text_in_r[16]$_DFFE_PP_  (.D(_00524_),
    .CK(clknet_leaf_0_clk),
    .Q(\text_in_r[16] ),
    .QN(_00462_));
 DFF_X2 \text_in_r[17]$_DFFE_PP_  (.D(_00525_),
    .CK(clknet_leaf_97_clk),
    .Q(\text_in_r[17] ),
    .QN(_00461_));
 DFF_X2 \text_in_r[18]$_DFFE_PP_  (.D(_00526_),
    .CK(clknet_leaf_97_clk),
    .Q(\text_in_r[18] ),
    .QN(_00463_));
 DFF_X1 \text_in_r[19]$_DFFE_PP_  (.D(_00527_),
    .CK(clknet_leaf_97_clk),
    .Q(\text_in_r[19] ),
    .QN(_14236_));
 DFF_X2 \text_in_r[1]$_DFFE_PP_  (.D(_00528_),
    .CK(clknet_leaf_19_clk),
    .Q(\text_in_r[1] ),
    .QN(_00405_));
 DFF_X2 \text_in_r[20]$_DFFE_PP_  (.D(_00529_),
    .CK(clknet_leaf_97_clk),
    .Q(\text_in_r[20] ),
    .QN(_14235_));
 DFF_X2 \text_in_r[21]$_DFFE_PP_  (.D(_00530_),
    .CK(clknet_leaf_0_clk),
    .Q(\text_in_r[21] ),
    .QN(_14234_));
 DFF_X1 \text_in_r[22]$_DFFE_PP_  (.D(_00531_),
    .CK(clknet_leaf_20_clk),
    .Q(\text_in_r[22] ),
    .QN(_14233_));
 DFF_X1 \text_in_r[23]$_DFFE_PP_  (.D(_00532_),
    .CK(clknet_leaf_20_clk),
    .Q(\text_in_r[23] ),
    .QN(_14232_));
 DFF_X1 \text_in_r[24]$_DFFE_PP_  (.D(_00533_),
    .CK(clknet_leaf_12_clk),
    .Q(\text_in_r[24] ),
    .QN(_00450_));
 DFF_X2 \text_in_r[25]$_DFFE_PP_  (.D(_00534_),
    .CK(clknet_leaf_17_clk),
    .Q(\text_in_r[25] ),
    .QN(_00449_));
 DFF_X1 \text_in_r[26]$_DFFE_PP_  (.D(_00535_),
    .CK(clknet_leaf_13_clk),
    .Q(\text_in_r[26] ),
    .QN(_00451_));
 DFF_X2 \text_in_r[27]$_DFFE_PP_  (.D(_00536_),
    .CK(clknet_leaf_13_clk),
    .Q(\text_in_r[27] ),
    .QN(_14231_));
 DFF_X2 \text_in_r[28]$_DFFE_PP_  (.D(_00537_),
    .CK(clknet_leaf_17_clk),
    .Q(\text_in_r[28] ),
    .QN(_14230_));
 DFF_X1 \text_in_r[29]$_DFFE_PP_  (.D(_00538_),
    .CK(clknet_leaf_4_clk),
    .Q(\text_in_r[29] ),
    .QN(_14229_));
 DFF_X1 \text_in_r[2]$_DFFE_PP_  (.D(_00539_),
    .CK(clknet_leaf_10_clk),
    .Q(\text_in_r[2] ),
    .QN(_00407_));
 DFF_X2 \text_in_r[30]$_DFFE_PP_  (.D(_00540_),
    .CK(clknet_leaf_13_clk),
    .Q(\text_in_r[30] ),
    .QN(_14228_));
 DFF_X1 \text_in_r[31]$_DFFE_PP_  (.D(_00541_),
    .CK(clknet_leaf_13_clk),
    .Q(\text_in_r[31] ),
    .QN(_14227_));
 DFF_X1 \text_in_r[32]$_DFFE_PP_  (.D(_00542_),
    .CK(clknet_leaf_57_clk),
    .Q(\text_in_r[32] ),
    .QN(_00483_));
 DFF_X1 \text_in_r[33]$_DFFE_PP_  (.D(_00543_),
    .CK(clknet_leaf_52_clk),
    .Q(\text_in_r[33] ),
    .QN(_00482_));
 DFF_X1 \text_in_r[34]$_DFFE_PP_  (.D(_00544_),
    .CK(clknet_leaf_51_clk),
    .Q(\text_in_r[34] ),
    .QN(_00484_));
 DFF_X1 \text_in_r[35]$_DFFE_PP_  (.D(_00545_),
    .CK(clknet_leaf_50_clk),
    .Q(\text_in_r[35] ),
    .QN(_14226_));
 DFF_X1 \text_in_r[36]$_DFFE_PP_  (.D(_00546_),
    .CK(clknet_leaf_48_clk),
    .Q(\text_in_r[36] ),
    .QN(_14225_));
 DFF_X1 \text_in_r[37]$_DFFE_PP_  (.D(_00547_),
    .CK(clknet_leaf_47_clk),
    .Q(\text_in_r[37] ),
    .QN(_14224_));
 DFF_X1 \text_in_r[38]$_DFFE_PP_  (.D(_00548_),
    .CK(clknet_leaf_52_clk),
    .Q(\text_in_r[38] ),
    .QN(_14223_));
 DFF_X1 \text_in_r[39]$_DFFE_PP_  (.D(_00549_),
    .CK(clknet_leaf_54_clk),
    .Q(\text_in_r[39] ),
    .QN(_14222_));
 DFF_X1 \text_in_r[3]$_DFFE_PP_  (.D(_00550_),
    .CK(clknet_leaf_15_clk),
    .Q(\text_in_r[3] ),
    .QN(_14221_));
 DFF_X1 \text_in_r[40]$_DFFE_PP_  (.D(_00551_),
    .CK(clknet_leaf_58_clk),
    .Q(\text_in_r[40] ),
    .QN(_00471_));
 DFF_X1 \text_in_r[41]$_DFFE_PP_  (.D(_00552_),
    .CK(clknet_leaf_58_clk),
    .Q(\text_in_r[41] ),
    .QN(_00470_));
 DFF_X1 \text_in_r[42]$_DFFE_PP_  (.D(_00553_),
    .CK(clknet_leaf_53_clk),
    .Q(\text_in_r[42] ),
    .QN(_00472_));
 DFF_X1 \text_in_r[43]$_DFFE_PP_  (.D(_00554_),
    .CK(clknet_leaf_70_clk),
    .Q(\text_in_r[43] ),
    .QN(_14220_));
 DFF_X1 \text_in_r[44]$_DFFE_PP_  (.D(_00555_),
    .CK(clknet_leaf_68_clk),
    .Q(\text_in_r[44] ),
    .QN(_14219_));
 DFF_X1 \text_in_r[45]$_DFFE_PP_  (.D(_00556_),
    .CK(clknet_leaf_59_clk),
    .Q(\text_in_r[45] ),
    .QN(_14218_));
 DFF_X1 \text_in_r[46]$_DFFE_PP_  (.D(_00557_),
    .CK(clknet_leaf_69_clk),
    .Q(\text_in_r[46] ),
    .QN(_14217_));
 DFF_X1 \text_in_r[47]$_DFFE_PP_  (.D(_00558_),
    .CK(clknet_leaf_69_clk),
    .Q(\text_in_r[47] ),
    .QN(_14216_));
 DFF_X1 \text_in_r[48]$_DFFE_PP_  (.D(_00559_),
    .CK(clknet_leaf_58_clk),
    .Q(\text_in_r[48] ),
    .QN(_00459_));
 DFF_X2 \text_in_r[49]$_DFFE_PP_  (.D(_00560_),
    .CK(clknet_leaf_60_clk),
    .Q(\text_in_r[49] ),
    .QN(_00458_));
 DFF_X1 \text_in_r[4]$_DFFE_PP_  (.D(_00561_),
    .CK(clknet_leaf_11_clk),
    .Q(\text_in_r[4] ),
    .QN(_14215_));
 DFF_X1 \text_in_r[50]$_DFFE_PP_  (.D(_00562_),
    .CK(clknet_leaf_61_clk),
    .Q(\text_in_r[50] ),
    .QN(_00460_));
 DFF_X1 \text_in_r[51]$_DFFE_PP_  (.D(_00563_),
    .CK(clknet_leaf_58_clk),
    .Q(\text_in_r[51] ),
    .QN(_14214_));
 DFF_X1 \text_in_r[52]$_DFFE_PP_  (.D(_00564_),
    .CK(clknet_leaf_60_clk),
    .Q(\text_in_r[52] ),
    .QN(_14213_));
 DFF_X1 \text_in_r[53]$_DFFE_PP_  (.D(_00565_),
    .CK(clknet_leaf_59_clk),
    .Q(\text_in_r[53] ),
    .QN(_14212_));
 DFF_X1 \text_in_r[54]$_DFFE_PP_  (.D(_00566_),
    .CK(clknet_leaf_68_clk),
    .Q(\text_in_r[54] ),
    .QN(_14211_));
 DFF_X1 \text_in_r[55]$_DFFE_PP_  (.D(_00567_),
    .CK(clknet_leaf_61_clk),
    .Q(\text_in_r[55] ),
    .QN(_14210_));
 DFF_X1 \text_in_r[56]$_DFFE_PP_  (.D(_00568_),
    .CK(clknet_leaf_62_clk),
    .Q(\text_in_r[56] ),
    .QN(_00447_));
 DFF_X2 \text_in_r[57]$_DFFE_PP_  (.D(_00569_),
    .CK(clknet_leaf_61_clk),
    .Q(\text_in_r[57] ),
    .QN(_00446_));
 DFF_X1 \text_in_r[58]$_DFFE_PP_  (.D(_00570_),
    .CK(clknet_leaf_62_clk),
    .Q(\text_in_r[58] ),
    .QN(_00448_));
 DFF_X1 \text_in_r[59]$_DFFE_PP_  (.D(_00571_),
    .CK(clknet_leaf_61_clk),
    .Q(\text_in_r[59] ),
    .QN(_14209_));
 DFF_X1 \text_in_r[5]$_DFFE_PP_  (.D(_00572_),
    .CK(clknet_leaf_12_clk),
    .Q(\text_in_r[5] ),
    .QN(_14208_));
 DFF_X1 \text_in_r[60]$_DFFE_PP_  (.D(_00573_),
    .CK(clknet_leaf_61_clk),
    .Q(\text_in_r[60] ),
    .QN(_14207_));
 DFF_X1 \text_in_r[61]$_DFFE_PP_  (.D(_00574_),
    .CK(clknet_leaf_60_clk),
    .Q(\text_in_r[61] ),
    .QN(_14206_));
 DFF_X1 \text_in_r[62]$_DFFE_PP_  (.D(_00575_),
    .CK(clknet_leaf_61_clk),
    .Q(\text_in_r[62] ),
    .QN(_14205_));
 DFF_X1 \text_in_r[63]$_DFFE_PP_  (.D(_00576_),
    .CK(clknet_leaf_61_clk),
    .Q(\text_in_r[63] ),
    .QN(_14204_));
 DFF_X1 \text_in_r[64]$_DFFE_PP_  (.D(_00577_),
    .CK(clknet_leaf_52_clk),
    .Q(\text_in_r[64] ),
    .QN(_00480_));
 DFF_X1 \text_in_r[65]$_DFFE_PP_  (.D(_00578_),
    .CK(clknet_leaf_39_clk),
    .Q(\text_in_r[65] ),
    .QN(_00479_));
 DFF_X1 \text_in_r[66]$_DFFE_PP_  (.D(_00579_),
    .CK(clknet_leaf_46_clk),
    .Q(\text_in_r[66] ),
    .QN(_00481_));
 DFF_X2 \text_in_r[67]$_DFFE_PP_  (.D(_00580_),
    .CK(clknet_leaf_49_clk),
    .Q(\text_in_r[67] ),
    .QN(_14203_));
 DFF_X1 \text_in_r[68]$_DFFE_PP_  (.D(_00581_),
    .CK(clknet_leaf_50_clk),
    .Q(\text_in_r[68] ),
    .QN(_14202_));
 DFF_X2 \text_in_r[69]$_DFFE_PP_  (.D(_00582_),
    .CK(clknet_leaf_48_clk),
    .Q(\text_in_r[69] ),
    .QN(_14201_));
 DFF_X1 \text_in_r[6]$_DFFE_PP_  (.D(_00583_),
    .CK(clknet_leaf_9_clk),
    .Q(\text_in_r[6] ),
    .QN(_14200_));
 DFF_X1 \text_in_r[70]$_DFFE_PP_  (.D(_00584_),
    .CK(clknet_leaf_46_clk),
    .Q(\text_in_r[70] ),
    .QN(_14199_));
 DFF_X1 \text_in_r[71]$_DFFE_PP_  (.D(_00585_),
    .CK(clknet_leaf_46_clk),
    .Q(\text_in_r[71] ),
    .QN(_14198_));
 DFF_X1 \text_in_r[72]$_DFFE_PP_  (.D(_00586_),
    .CK(clknet_leaf_55_clk),
    .Q(\text_in_r[72] ),
    .QN(_00468_));
 DFF_X2 \text_in_r[73]$_DFFE_PP_  (.D(_00587_),
    .CK(clknet_leaf_27_clk),
    .Q(\text_in_r[73] ),
    .QN(_00467_));
 DFF_X1 \text_in_r[74]$_DFFE_PP_  (.D(_00588_),
    .CK(clknet_leaf_55_clk),
    .Q(\text_in_r[74] ),
    .QN(_00469_));
 DFF_X2 \text_in_r[75]$_DFFE_PP_  (.D(_00589_),
    .CK(clknet_leaf_51_clk),
    .Q(\text_in_r[75] ),
    .QN(_14197_));
 DFF_X2 \text_in_r[76]$_DFFE_PP_  (.D(_00590_),
    .CK(clknet_leaf_31_clk),
    .Q(\text_in_r[76] ),
    .QN(_14196_));
 DFF_X2 \text_in_r[77]$_DFFE_PP_  (.D(_00591_),
    .CK(clknet_leaf_56_clk),
    .Q(\text_in_r[77] ),
    .QN(_14195_));
 DFF_X1 \text_in_r[78]$_DFFE_PP_  (.D(_00592_),
    .CK(clknet_leaf_8_clk),
    .Q(\text_in_r[78] ),
    .QN(_14194_));
 DFF_X1 \text_in_r[79]$_DFFE_PP_  (.D(_00593_),
    .CK(clknet_leaf_53_clk),
    .Q(\text_in_r[79] ),
    .QN(_14193_));
 DFF_X1 \text_in_r[7]$_DFFE_PP_  (.D(_00594_),
    .CK(clknet_leaf_11_clk),
    .Q(\text_in_r[7] ),
    .QN(_14192_));
 DFF_X1 \text_in_r[80]$_DFFE_PP_  (.D(_00595_),
    .CK(clknet_leaf_54_clk),
    .Q(\text_in_r[80] ),
    .QN(_00456_));
 DFF_X2 \text_in_r[81]$_DFFE_PP_  (.D(_00596_),
    .CK(clknet_leaf_54_clk),
    .Q(\text_in_r[81] ),
    .QN(_00455_));
 DFF_X1 \text_in_r[82]$_DFFE_PP_  (.D(_00597_),
    .CK(clknet_leaf_55_clk),
    .Q(\text_in_r[82] ),
    .QN(_00457_));
 DFF_X1 \text_in_r[83]$_DFFE_PP_  (.D(_00598_),
    .CK(clknet_leaf_54_clk),
    .Q(\text_in_r[83] ),
    .QN(_14191_));
 DFF_X2 \text_in_r[84]$_DFFE_PP_  (.D(_00599_),
    .CK(clknet_leaf_57_clk),
    .Q(\text_in_r[84] ),
    .QN(_14190_));
 DFF_X1 \text_in_r[85]$_DFFE_PP_  (.D(_00600_),
    .CK(clknet_leaf_62_clk),
    .Q(\text_in_r[85] ),
    .QN(_14189_));
 DFF_X1 \text_in_r[86]$_DFFE_PP_  (.D(_00601_),
    .CK(clknet_leaf_53_clk),
    .Q(\text_in_r[86] ),
    .QN(_14188_));
 DFF_X1 \text_in_r[87]$_DFFE_PP_  (.D(_00602_),
    .CK(clknet_leaf_53_clk),
    .Q(\text_in_r[87] ),
    .QN(_14187_));
 DFF_X1 \text_in_r[88]$_DFFE_PP_  (.D(_00603_),
    .CK(clknet_leaf_47_clk),
    .Q(\text_in_r[88] ),
    .QN(_00444_));
 DFF_X1 \text_in_r[89]$_DFFE_PP_  (.D(_00604_),
    .CK(clknet_leaf_48_clk),
    .Q(\text_in_r[89] ),
    .QN(_00443_));
 DFF_X1 \text_in_r[8]$_DFFE_PP_  (.D(_00605_),
    .CK(clknet_leaf_30_clk),
    .Q(\text_in_r[8] ),
    .QN(_00474_));
 DFF_X1 \text_in_r[90]$_DFFE_PP_  (.D(_00606_),
    .CK(clknet_leaf_52_clk),
    .Q(\text_in_r[90] ),
    .QN(_00445_));
 DFF_X1 \text_in_r[91]$_DFFE_PP_  (.D(_00607_),
    .CK(clknet_leaf_48_clk),
    .Q(\text_in_r[91] ),
    .QN(_14186_));
 DFF_X2 \text_in_r[92]$_DFFE_PP_  (.D(_00608_),
    .CK(clknet_leaf_49_clk),
    .Q(\text_in_r[92] ),
    .QN(_14185_));
 DFF_X1 \text_in_r[93]$_DFFE_PP_  (.D(_00609_),
    .CK(clknet_leaf_45_clk),
    .Q(\text_in_r[93] ),
    .QN(_14184_));
 DFF_X1 \text_in_r[94]$_DFFE_PP_  (.D(_00610_),
    .CK(clknet_leaf_46_clk),
    .Q(\text_in_r[94] ),
    .QN(_14183_));
 DFF_X1 \text_in_r[95]$_DFFE_PP_  (.D(_00611_),
    .CK(clknet_leaf_46_clk),
    .Q(\text_in_r[95] ),
    .QN(_14182_));
 DFF_X1 \text_in_r[96]$_DFFE_PP_  (.D(_00612_),
    .CK(clknet_leaf_30_clk),
    .Q(\text_in_r[96] ),
    .QN(_00477_));
 DFF_X1 \text_in_r[97]$_DFFE_PP_  (.D(_00613_),
    .CK(clknet_leaf_36_clk),
    .Q(\text_in_r[97] ),
    .QN(_00476_));
 DFF_X1 \text_in_r[98]$_DFFE_PP_  (.D(_00614_),
    .CK(clknet_leaf_28_clk),
    .Q(\text_in_r[98] ),
    .QN(_00478_));
 DFF_X1 \text_in_r[99]$_DFFE_PP_  (.D(_00615_),
    .CK(clknet_leaf_32_clk),
    .Q(\text_in_r[99] ),
    .QN(_14181_));
 DFF_X1 \text_in_r[9]$_DFFE_PP_  (.D(_00616_),
    .CK(clknet_leaf_5_clk),
    .Q(\text_in_r[9] ),
    .QN(_00473_));
 DFF_X2 \text_out[0]$_DFF_P_  (.D(_00265_),
    .CK(clknet_leaf_14_clk),
    .Q(net357),
    .QN(_14395_));
 DFF_X1 \text_out[100]$_DFF_P_  (.D(_00165_),
    .CK(clknet_leaf_34_clk),
    .Q(net358),
    .QN(_14396_));
 DFF_X2 \text_out[101]$_DFF_P_  (.D(_00166_),
    .CK(clknet_leaf_51_clk),
    .Q(net359),
    .QN(_14397_));
 DFF_X2 \text_out[102]$_DFF_P_  (.D(_00167_),
    .CK(clknet_leaf_41_clk),
    .Q(net360),
    .QN(_14398_));
 DFF_X1 \text_out[103]$_DFF_P_  (.D(_00168_),
    .CK(clknet_leaf_38_clk),
    .Q(net361),
    .QN(_14399_));
 DFF_X1 \text_out[104]$_DFF_P_  (.D(_00169_),
    .CK(clknet_leaf_94_clk),
    .Q(net362),
    .QN(_14400_));
 DFF_X1 \text_out[105]$_DFF_P_  (.D(_00170_),
    .CK(clknet_leaf_28_clk),
    .Q(net363),
    .QN(_14401_));
 DFF_X2 \text_out[106]$_DFF_P_  (.D(_00171_),
    .CK(clknet_leaf_58_clk),
    .Q(net364),
    .QN(_14402_));
 DFF_X1 \text_out[107]$_DFF_P_  (.D(_00172_),
    .CK(clknet_leaf_73_clk),
    .Q(net365),
    .QN(_14403_));
 DFF_X1 \text_out[108]$_DFF_P_  (.D(_00173_),
    .CK(clknet_leaf_73_clk),
    .Q(net366),
    .QN(_14404_));
 DFF_X1 \text_out[109]$_DFF_P_  (.D(_00174_),
    .CK(clknet_leaf_91_clk),
    .Q(net367),
    .QN(_14405_));
 DFF_X1 \text_out[10]$_DFF_P_  (.D(_00195_),
    .CK(clknet_leaf_0_clk),
    .Q(net368),
    .QN(_14406_));
 DFF_X1 \text_out[110]$_DFF_P_  (.D(_00175_),
    .CK(clknet_leaf_94_clk),
    .Q(net369),
    .QN(_14407_));
 DFF_X1 \text_out[111]$_DFF_P_  (.D(_00176_),
    .CK(clknet_leaf_92_clk),
    .Q(net370),
    .QN(_14408_));
 DFF_X1 \text_out[112]$_DFF_P_  (.D(_00177_),
    .CK(clknet_leaf_93_clk),
    .Q(net371),
    .QN(_14409_));
 DFF_X1 \text_out[113]$_DFF_P_  (.D(_00178_),
    .CK(clknet_leaf_82_clk),
    .Q(net372),
    .QN(_14410_));
 DFF_X1 \text_out[114]$_DFF_P_  (.D(_00179_),
    .CK(clknet_leaf_92_clk),
    .Q(net373),
    .QN(_14411_));
 DFF_X1 \text_out[115]$_DFF_P_  (.D(_00180_),
    .CK(clknet_leaf_84_clk),
    .Q(net374),
    .QN(_14412_));
 DFF_X1 \text_out[116]$_DFF_P_  (.D(_00181_),
    .CK(clknet_leaf_85_clk),
    .Q(net375),
    .QN(_14413_));
 DFF_X1 \text_out[117]$_DFF_P_  (.D(_00182_),
    .CK(clknet_leaf_82_clk),
    .Q(net376),
    .QN(_14414_));
 DFF_X1 \text_out[118]$_DFF_P_  (.D(_00183_),
    .CK(clknet_leaf_86_clk),
    .Q(net377),
    .QN(_14415_));
 DFF_X1 \text_out[119]$_DFF_P_  (.D(_00184_),
    .CK(clknet_leaf_83_clk),
    .Q(net378),
    .QN(_14416_));
 DFF_X1 \text_out[11]$_DFF_P_  (.D(_00196_),
    .CK(clknet_leaf_0_clk),
    .Q(net379),
    .QN(_14417_));
 DFF_X1 \text_out[120]$_DFF_P_  (.D(_00185_),
    .CK(clknet_leaf_73_clk),
    .Q(net380),
    .QN(_14418_));
 DFF_X1 \text_out[121]$_DFF_P_  (.D(_00186_),
    .CK(clknet_leaf_94_clk),
    .Q(net381),
    .QN(_14419_));
 DFF_X1 \text_out[122]$_DFF_P_  (.D(_00187_),
    .CK(clknet_leaf_92_clk),
    .Q(net382),
    .QN(_14420_));
 DFF_X1 \text_out[123]$_DFF_P_  (.D(_00188_),
    .CK(clknet_leaf_94_clk),
    .Q(net383),
    .QN(_14421_));
 DFF_X1 \text_out[124]$_DFF_P_  (.D(_00189_),
    .CK(clknet_leaf_72_clk),
    .Q(net384),
    .QN(_14422_));
 DFF_X1 \text_out[125]$_DFF_P_  (.D(_00190_),
    .CK(clknet_leaf_93_clk),
    .Q(net385),
    .QN(_14423_));
 DFF_X1 \text_out[126]$_DFF_P_  (.D(_00191_),
    .CK(clknet_leaf_67_clk),
    .Q(net386),
    .QN(_14424_));
 DFF_X2 \text_out[127]$_DFF_P_  (.D(_00192_),
    .CK(clknet_leaf_76_clk),
    .Q(net387),
    .QN(_14425_));
 DFF_X1 \text_out[12]$_DFF_P_  (.D(_00197_),
    .CK(clknet_leaf_0_clk),
    .Q(net388),
    .QN(_14426_));
 DFF_X1 \text_out[13]$_DFF_P_  (.D(_00198_),
    .CK(clknet_leaf_0_clk),
    .Q(net389),
    .QN(_14427_));
 DFF_X1 \text_out[14]$_DFF_P_  (.D(_00199_),
    .CK(clknet_leaf_13_clk),
    .Q(net390),
    .QN(_14428_));
 DFF_X1 \text_out[15]$_DFF_P_  (.D(_00200_),
    .CK(clknet_leaf_20_clk),
    .Q(net391),
    .QN(_14429_));
 DFF_X2 \text_out[16]$_DFF_P_  (.D(_00201_),
    .CK(clknet_leaf_4_clk),
    .Q(net392),
    .QN(_14430_));
 DFF_X2 \text_out[17]$_DFF_P_  (.D(_00202_),
    .CK(clknet_leaf_88_clk),
    .Q(net393),
    .QN(_14431_));
 DFF_X1 \text_out[18]$_DFF_P_  (.D(_00203_),
    .CK(clknet_leaf_1_clk),
    .Q(net394),
    .QN(_14432_));
 DFF_X1 \text_out[19]$_DFF_P_  (.D(_00204_),
    .CK(clknet_leaf_97_clk),
    .Q(net395),
    .QN(_14433_));
 DFF_X2 \text_out[1]$_DFF_P_  (.D(_00266_),
    .CK(clknet_leaf_14_clk),
    .Q(net396),
    .QN(_14434_));
 DFF_X2 \text_out[20]$_DFF_P_  (.D(_00205_),
    .CK(clknet_leaf_88_clk),
    .Q(net397),
    .QN(_14435_));
 DFF_X1 \text_out[21]$_DFF_P_  (.D(_00206_),
    .CK(clknet_leaf_96_clk),
    .Q(net398),
    .QN(_14436_));
 DFF_X1 \text_out[22]$_DFF_P_  (.D(_00207_),
    .CK(clknet_leaf_2_clk),
    .Q(net399),
    .QN(_14437_));
 DFF_X2 \text_out[23]$_DFF_P_  (.D(_00208_),
    .CK(clknet_leaf_88_clk),
    .Q(net400),
    .QN(_14438_));
 DFF_X2 \text_out[24]$_DFF_P_  (.D(_00209_),
    .CK(clknet_leaf_11_clk),
    .Q(net401),
    .QN(_14439_));
 DFF_X2 \text_out[25]$_DFF_P_  (.D(_00210_),
    .CK(clknet_leaf_12_clk),
    .Q(net402),
    .QN(_14440_));
 DFF_X2 \text_out[26]$_DFF_P_  (.D(_00211_),
    .CK(clknet_leaf_10_clk),
    .Q(net403),
    .QN(_14441_));
 DFF_X2 \text_out[27]$_DFF_P_  (.D(_00212_),
    .CK(clknet_leaf_14_clk),
    .Q(net404),
    .QN(_14442_));
 DFF_X2 \text_out[28]$_DFF_P_  (.D(_00213_),
    .CK(clknet_leaf_4_clk),
    .Q(net405),
    .QN(_14443_));
 DFF_X1 \text_out[29]$_DFF_P_  (.D(_00214_),
    .CK(clknet_leaf_18_clk),
    .Q(net406),
    .QN(_14444_));
 DFF_X1 \text_out[2]$_DFF_P_  (.D(_00267_),
    .CK(clknet_leaf_19_clk),
    .Q(net407),
    .QN(_14445_));
 DFF_X1 \text_out[30]$_DFF_P_  (.D(_00215_),
    .CK(clknet_leaf_13_clk),
    .Q(net408),
    .QN(_14446_));
 DFF_X1 \text_out[31]$_DFF_P_  (.D(_00216_),
    .CK(clknet_leaf_18_clk),
    .Q(net409),
    .QN(_14447_));
 DFF_X1 \text_out[32]$_DFF_P_  (.D(_00217_),
    .CK(clknet_leaf_47_clk),
    .Q(net410),
    .QN(_14448_));
 DFF_X2 \text_out[33]$_DFF_P_  (.D(_00218_),
    .CK(clknet_leaf_52_clk),
    .Q(net411),
    .QN(_14449_));
 DFF_X2 \text_out[34]$_DFF_P_  (.D(_00219_),
    .CK(clknet_leaf_39_clk),
    .Q(net412),
    .QN(_14450_));
 DFF_X1 \text_out[35]$_DFF_P_  (.D(_00220_),
    .CK(clknet_leaf_43_clk),
    .Q(net413),
    .QN(_14451_));
 DFF_X1 \text_out[36]$_DFF_P_  (.D(_00221_),
    .CK(clknet_leaf_49_clk),
    .Q(net414),
    .QN(_14452_));
 DFF_X1 \text_out[37]$_DFF_P_  (.D(_00222_),
    .CK(clknet_leaf_49_clk),
    .Q(net415),
    .QN(_14453_));
 DFF_X1 \text_out[38]$_DFF_P_  (.D(_00223_),
    .CK(clknet_leaf_50_clk),
    .Q(net416),
    .QN(_14454_));
 DFF_X2 \text_out[39]$_DFF_P_  (.D(_00224_),
    .CK(clknet_leaf_50_clk),
    .Q(net417),
    .QN(_14455_));
 DFF_X1 \text_out[3]$_DFF_P_  (.D(_00268_),
    .CK(clknet_leaf_21_clk),
    .Q(net418),
    .QN(_14456_));
 DFF_X1 \text_out[40]$_DFF_P_  (.D(_00225_),
    .CK(clknet_leaf_71_clk),
    .Q(net419),
    .QN(_14457_));
 DFF_X2 \text_out[41]$_DFF_P_  (.D(_00226_),
    .CK(clknet_leaf_60_clk),
    .Q(net420),
    .QN(_14458_));
 DFF_X1 \text_out[42]$_DFF_P_  (.D(_00227_),
    .CK(clknet_leaf_65_clk),
    .Q(net421),
    .QN(_14459_));
 DFF_X1 \text_out[43]$_DFF_P_  (.D(_00228_),
    .CK(clknet_leaf_59_clk),
    .Q(net422),
    .QN(_14460_));
 DFF_X1 \text_out[44]$_DFF_P_  (.D(_00229_),
    .CK(clknet_leaf_59_clk),
    .Q(net423),
    .QN(_14461_));
 DFF_X1 \text_out[45]$_DFF_P_  (.D(_00230_),
    .CK(clknet_leaf_60_clk),
    .Q(net424),
    .QN(_14462_));
 DFF_X2 \text_out[46]$_DFF_P_  (.D(_00231_),
    .CK(clknet_leaf_69_clk),
    .Q(net425),
    .QN(_14463_));
 DFF_X2 \text_out[47]$_DFF_P_  (.D(_00232_),
    .CK(clknet_leaf_70_clk),
    .Q(net426),
    .QN(_14464_));
 DFF_X1 \text_out[48]$_DFF_P_  (.D(_00233_),
    .CK(clknet_leaf_94_clk),
    .Q(net427),
    .QN(_14465_));
 DFF_X2 \text_out[49]$_DFF_P_  (.D(_00234_),
    .CK(clknet_leaf_82_clk),
    .Q(net428),
    .QN(_14466_));
 DFF_X1 \text_out[4]$_DFF_P_  (.D(_00269_),
    .CK(clknet_leaf_22_clk),
    .Q(net429),
    .QN(_14467_));
 DFF_X1 \text_out[50]$_DFF_P_  (.D(_00235_),
    .CK(clknet_leaf_65_clk),
    .Q(net430),
    .QN(_14468_));
 DFF_X1 \text_out[51]$_DFF_P_  (.D(_00236_),
    .CK(clknet_leaf_58_clk),
    .Q(net431),
    .QN(_14469_));
 DFF_X1 \text_out[52]$_DFF_P_  (.D(_00237_),
    .CK(clknet_leaf_93_clk),
    .Q(net432),
    .QN(_14470_));
 DFF_X1 \text_out[53]$_DFF_P_  (.D(_00238_),
    .CK(clknet_leaf_84_clk),
    .Q(net433),
    .QN(_14471_));
 DFF_X1 \text_out[54]$_DFF_P_  (.D(_00239_),
    .CK(clknet_leaf_86_clk),
    .Q(net434),
    .QN(_14472_));
 DFF_X1 \text_out[55]$_DFF_P_  (.D(_00240_),
    .CK(clknet_leaf_60_clk),
    .Q(net435),
    .QN(_14473_));
 DFF_X1 \text_out[56]$_DFF_P_  (.D(_00241_),
    .CK(clknet_leaf_65_clk),
    .Q(net436),
    .QN(_14474_));
 DFF_X1 \text_out[57]$_DFF_P_  (.D(_00242_),
    .CK(clknet_leaf_65_clk),
    .Q(net437),
    .QN(_14475_));
 DFF_X1 \text_out[58]$_DFF_P_  (.D(_00243_),
    .CK(clknet_leaf_65_clk),
    .Q(net438),
    .QN(_14476_));
 DFF_X1 \text_out[59]$_DFF_P_  (.D(_00244_),
    .CK(clknet_leaf_68_clk),
    .Q(net439),
    .QN(_14477_));
 DFF_X2 \text_out[5]$_DFF_P_  (.D(_00270_),
    .CK(clknet_leaf_11_clk),
    .Q(net440),
    .QN(_14478_));
 DFF_X1 \text_out[60]$_DFF_P_  (.D(_00245_),
    .CK(clknet_leaf_68_clk),
    .Q(net441),
    .QN(_14479_));
 DFF_X1 \text_out[61]$_DFF_P_  (.D(_00246_),
    .CK(clknet_leaf_66_clk),
    .Q(net442),
    .QN(_14480_));
 DFF_X1 \text_out[62]$_DFF_P_  (.D(_00247_),
    .CK(clknet_leaf_64_clk),
    .Q(net443),
    .QN(_14481_));
 DFF_X1 \text_out[63]$_DFF_P_  (.D(_00248_),
    .CK(clknet_leaf_65_clk),
    .Q(net444),
    .QN(_14482_));
 DFF_X1 \text_out[64]$_DFF_P_  (.D(_00249_),
    .CK(clknet_leaf_52_clk),
    .Q(net445),
    .QN(_14483_));
 DFF_X1 \text_out[65]$_DFF_P_  (.D(_00250_),
    .CK(clknet_leaf_39_clk),
    .Q(net446),
    .QN(_14484_));
 DFF_X1 \text_out[66]$_DFF_P_  (.D(_00251_),
    .CK(clknet_leaf_39_clk),
    .Q(net447),
    .QN(_14485_));
 DFF_X1 \text_out[67]$_DFF_P_  (.D(_00252_),
    .CK(clknet_leaf_41_clk),
    .Q(net448),
    .QN(_14486_));
 DFF_X1 \text_out[68]$_DFF_P_  (.D(_00253_),
    .CK(clknet_leaf_41_clk),
    .Q(net449),
    .QN(_14487_));
 DFF_X1 \text_out[69]$_DFF_P_  (.D(_00254_),
    .CK(clknet_leaf_49_clk),
    .Q(net450),
    .QN(_14488_));
 DFF_X1 \text_out[6]$_DFF_P_  (.D(_00271_),
    .CK(clknet_leaf_22_clk),
    .Q(net451),
    .QN(_14489_));
 DFF_X2 \text_out[70]$_DFF_P_  (.D(_00255_),
    .CK(clknet_leaf_41_clk),
    .Q(net452),
    .QN(_14490_));
 DFF_X1 \text_out[71]$_DFF_P_  (.D(_00256_),
    .CK(clknet_leaf_48_clk),
    .Q(net453),
    .QN(_14491_));
 DFF_X2 \text_out[72]$_DFF_P_  (.D(_00257_),
    .CK(clknet_leaf_56_clk),
    .Q(net454),
    .QN(_14492_));
 DFF_X1 \text_out[73]$_DFF_P_  (.D(_00258_),
    .CK(clknet_leaf_22_clk),
    .Q(net455),
    .QN(_14493_));
 DFF_X2 \text_out[74]$_DFF_P_  (.D(_00259_),
    .CK(clknet_leaf_55_clk),
    .Q(net456),
    .QN(_14494_));
 DFF_X2 \text_out[75]$_DFF_P_  (.D(_00260_),
    .CK(clknet_leaf_55_clk),
    .Q(net457),
    .QN(_14495_));
 DFF_X2 \text_out[76]$_DFF_P_  (.D(_00261_),
    .CK(clknet_leaf_56_clk),
    .Q(net458),
    .QN(_14496_));
 DFF_X1 \text_out[77]$_DFF_P_  (.D(_00262_),
    .CK(clknet_leaf_22_clk),
    .Q(net459),
    .QN(_14497_));
 DFF_X2 \text_out[78]$_DFF_P_  (.D(_00263_),
    .CK(clknet_leaf_79_clk),
    .Q(net460),
    .QN(_14498_));
 DFF_X1 \text_out[79]$_DFF_P_  (.D(_00264_),
    .CK(clknet_leaf_37_clk),
    .Q(net461),
    .QN(_14499_));
 DFF_X2 \text_out[7]$_DFF_P_  (.D(_00272_),
    .CK(clknet_leaf_14_clk),
    .Q(net462),
    .QN(_14500_));
 DFF_X1 \text_out[80]$_DFF_P_  (.D(_00273_),
    .CK(clknet_leaf_45_clk),
    .Q(net463),
    .QN(_14501_));
 DFF_X2 \text_out[81]$_DFF_P_  (.D(_00274_),
    .CK(clknet_leaf_54_clk),
    .Q(net464),
    .QN(_14502_));
 DFF_X2 \text_out[82]$_DFF_P_  (.D(_00275_),
    .CK(clknet_leaf_55_clk),
    .Q(net465),
    .QN(_14503_));
 DFF_X1 \text_out[83]$_DFF_P_  (.D(_00276_),
    .CK(clknet_leaf_53_clk),
    .Q(net466),
    .QN(_14504_));
 DFF_X1 \text_out[84]$_DFF_P_  (.D(_00277_),
    .CK(clknet_leaf_62_clk),
    .Q(net467),
    .QN(_14505_));
 DFF_X1 \text_out[85]$_DFF_P_  (.D(_00278_),
    .CK(clknet_leaf_44_clk),
    .Q(net468),
    .QN(_14506_));
 DFF_X1 \text_out[86]$_DFF_P_  (.D(_00279_),
    .CK(clknet_leaf_57_clk),
    .Q(net469),
    .QN(_14507_));
 DFF_X1 \text_out[87]$_DFF_P_  (.D(_00280_),
    .CK(clknet_leaf_67_clk),
    .Q(net470),
    .QN(_14508_));
 DFF_X1 \text_out[88]$_DFF_P_  (.D(_00281_),
    .CK(clknet_leaf_47_clk),
    .Q(net471),
    .QN(_14509_));
 DFF_X1 \text_out[89]$_DFF_P_  (.D(_00282_),
    .CK(clknet_leaf_45_clk),
    .Q(net472),
    .QN(_14510_));
 DFF_X1 \text_out[8]$_DFF_P_  (.D(_00193_),
    .CK(clknet_leaf_20_clk),
    .Q(net473),
    .QN(_14511_));
 DFF_X1 \text_out[90]$_DFF_P_  (.D(_00283_),
    .CK(clknet_leaf_53_clk),
    .Q(net474),
    .QN(_14512_));
 DFF_X1 \text_out[91]$_DFF_P_  (.D(_00284_),
    .CK(clknet_leaf_48_clk),
    .Q(net475),
    .QN(_14513_));
 DFF_X1 \text_out[92]$_DFF_P_  (.D(_00285_),
    .CK(clknet_leaf_45_clk),
    .Q(net476),
    .QN(_14514_));
 DFF_X1 \text_out[93]$_DFF_P_  (.D(_00286_),
    .CK(clknet_leaf_44_clk),
    .Q(net477),
    .QN(_14515_));
 DFF_X1 \text_out[94]$_DFF_P_  (.D(_00287_),
    .CK(clknet_leaf_45_clk),
    .Q(net478),
    .QN(_14516_));
 DFF_X1 \text_out[95]$_DFF_P_  (.D(_00288_),
    .CK(clknet_leaf_45_clk),
    .Q(net479),
    .QN(_14517_));
 DFF_X1 \text_out[96]$_DFF_P_  (.D(_00161_),
    .CK(clknet_leaf_31_clk),
    .Q(net480),
    .QN(_14518_));
 DFF_X2 \text_out[97]$_DFF_P_  (.D(_00162_),
    .CK(clknet_leaf_23_clk),
    .Q(net481),
    .QN(_14519_));
 DFF_X1 \text_out[98]$_DFF_P_  (.D(_00163_),
    .CK(clknet_leaf_37_clk),
    .Q(net482),
    .QN(_14520_));
 DFF_X1 \text_out[99]$_DFF_P_  (.D(_00164_),
    .CK(clknet_leaf_35_clk),
    .Q(net483),
    .QN(_14521_));
 DFF_X1 \text_out[9]$_DFF_P_  (.D(_00194_),
    .CK(clknet_leaf_0_clk),
    .Q(net484),
    .QN(_14180_));
 DFF_X1 \u0.r0.out[24]$_SDFF_PP1_  (.D(_00617_),
    .CK(clknet_leaf_9_clk),
    .Q(\u0.r0.out[24] ),
    .QN(_00432_));
 DFF_X1 \u0.r0.out[25]$_SDFF_PP0_  (.D(_00618_),
    .CK(clknet_leaf_12_clk),
    .Q(\u0.r0.out[25] ),
    .QN(_00433_));
 DFF_X1 \u0.r0.out[26]$_SDFF_PP0_  (.D(_00619_),
    .CK(clknet_leaf_7_clk),
    .Q(\u0.r0.out[26] ),
    .QN(_00434_));
 DFF_X1 \u0.r0.out[27]$_SDFF_PP0_  (.D(_00620_),
    .CK(clknet_leaf_5_clk),
    .Q(\u0.r0.out[27] ),
    .QN(_00435_));
 DFF_X1 \u0.r0.out[28]$_SDFF_PP0_  (.D(_00621_),
    .CK(clknet_leaf_7_clk),
    .Q(\u0.r0.out[28] ),
    .QN(_00436_));
 DFF_X1 \u0.r0.out[29]$_SDFF_PP0_  (.D(_00622_),
    .CK(clknet_leaf_7_clk),
    .Q(\u0.r0.out[29] ),
    .QN(_00437_));
 DFF_X1 \u0.r0.out[30]$_SDFF_PP0_  (.D(_00623_),
    .CK(clknet_leaf_6_clk),
    .Q(\u0.r0.out[30] ),
    .QN(_00438_));
 DFF_X1 \u0.r0.out[31]$_SDFF_PP0_  (.D(_00624_),
    .CK(clknet_leaf_9_clk),
    .Q(\u0.r0.out[31] ),
    .QN(_00439_));
 DFF_X2 \u0.r0.rcnt[0]$_SDFF_PP0_  (.D(_00625_),
    .CK(clknet_leaf_5_clk),
    .Q(\u0.r0.rcnt[0] ),
    .QN(\u0.r0.rcnt_next[0] ));
 DFF_X2 \u0.r0.rcnt[1]$_SDFF_PP0_  (.D(_00626_),
    .CK(clknet_leaf_5_clk),
    .Q(\u0.r0.rcnt[1] ),
    .QN(_15322_));
 DFF_X2 \u0.r0.rcnt[2]$_SDFF_PP0_  (.D(_00627_),
    .CK(clknet_leaf_12_clk),
    .Q(\u0.r0.rcnt[2] ),
    .QN(_14179_));
 DFF_X1 \u0.r0.rcnt[3]$_SDFF_PP0_  (.D(_00628_),
    .CK(clknet_leaf_5_clk),
    .Q(\u0.r0.rcnt[3] ),
    .QN(_14522_));
 DFF_X1 \u0.u0.d[0]$_DFF_P_  (.D(_00000_),
    .CK(clknet_leaf_85_clk),
    .Q(\u0.subword[24] ),
    .QN(_14523_));
 DFF_X2 \u0.u0.d[1]$_DFF_P_  (.D(_00001_),
    .CK(clknet_leaf_90_clk),
    .Q(\u0.subword[25] ),
    .QN(_14524_));
 DFF_X2 \u0.u0.d[2]$_DFF_P_  (.D(_00002_),
    .CK(clknet_leaf_90_clk),
    .Q(\u0.subword[26] ),
    .QN(_14525_));
 DFF_X2 \u0.u0.d[3]$_DFF_P_  (.D(_00003_),
    .CK(clknet_leaf_89_clk),
    .Q(\u0.subword[27] ),
    .QN(_14526_));
 DFF_X1 \u0.u0.d[4]$_DFF_P_  (.D(_00004_),
    .CK(clknet_leaf_90_clk),
    .Q(\u0.subword[28] ),
    .QN(_14527_));
 DFF_X1 \u0.u0.d[5]$_DFF_P_  (.D(_00005_),
    .CK(clknet_leaf_90_clk),
    .Q(\u0.subword[29] ),
    .QN(_14528_));
 DFF_X1 \u0.u0.d[6]$_DFF_P_  (.D(_00006_),
    .CK(clknet_leaf_89_clk),
    .Q(\u0.subword[30] ),
    .QN(_14529_));
 DFF_X1 \u0.u0.d[7]$_DFF_P_  (.D(_00007_),
    .CK(clknet_leaf_91_clk),
    .Q(\u0.subword[31] ),
    .QN(_14530_));
 DFF_X1 \u0.u1.d[0]$_DFF_P_  (.D(_00008_),
    .CK(clknet_leaf_6_clk),
    .Q(\u0.subword[16] ),
    .QN(_00425_));
 DFF_X1 \u0.u1.d[1]$_DFF_P_  (.D(_00009_),
    .CK(clknet_leaf_87_clk),
    .Q(\u0.subword[17] ),
    .QN(_00426_));
 DFF_X1 \u0.u1.d[2]$_DFF_P_  (.D(_00010_),
    .CK(clknet_leaf_87_clk),
    .Q(\u0.subword[18] ),
    .QN(_00408_));
 DFF_X1 \u0.u1.d[3]$_DFF_P_  (.D(_00011_),
    .CK(clknet_leaf_87_clk),
    .Q(\u0.subword[19] ),
    .QN(_00427_));
 DFF_X1 \u0.u1.d[4]$_DFF_P_  (.D(_00012_),
    .CK(clknet_leaf_85_clk),
    .Q(\u0.subword[20] ),
    .QN(_00428_));
 DFF_X1 \u0.u1.d[5]$_DFF_P_  (.D(_00013_),
    .CK(clknet_leaf_90_clk),
    .Q(\u0.subword[21] ),
    .QN(_00429_));
 DFF_X2 \u0.u1.d[6]$_DFF_P_  (.D(_00014_),
    .CK(clknet_leaf_3_clk),
    .Q(\u0.subword[22] ),
    .QN(_00430_));
 DFF_X1 \u0.u1.d[7]$_DFF_P_  (.D(_00015_),
    .CK(clknet_leaf_84_clk),
    .Q(\u0.subword[23] ),
    .QN(_00431_));
 DFF_X2 \u0.u2.d[0]$_DFF_P_  (.D(_00016_),
    .CK(clknet_leaf_24_clk),
    .Q(\u0.subword[8] ),
    .QN(_00418_));
 DFF_X2 \u0.u2.d[1]$_DFF_P_  (.D(_00017_),
    .CK(clknet_leaf_27_clk),
    .Q(\u0.subword[9] ),
    .QN(_00419_));
 DFF_X2 \u0.u2.d[2]$_DFF_P_  (.D(_00018_),
    .CK(clknet_leaf_24_clk),
    .Q(\u0.subword[10] ),
    .QN(_00410_));
 DFF_X1 \u0.u2.d[3]$_DFF_P_  (.D(_00019_),
    .CK(clknet_leaf_80_clk),
    .Q(\u0.subword[11] ),
    .QN(_00420_));
 DFF_X1 \u0.u2.d[4]$_DFF_P_  (.D(_00020_),
    .CK(clknet_leaf_8_clk),
    .Q(\u0.subword[12] ),
    .QN(_00421_));
 DFF_X1 \u0.u2.d[5]$_DFF_P_  (.D(_00021_),
    .CK(clknet_leaf_81_clk),
    .Q(\u0.subword[13] ),
    .QN(_00422_));
 DFF_X1 \u0.u2.d[6]$_DFF_P_  (.D(_00022_),
    .CK(clknet_leaf_7_clk),
    .Q(\u0.subword[14] ),
    .QN(_00423_));
 DFF_X1 \u0.u2.d[7]$_DFF_P_  (.D(_00023_),
    .CK(clknet_leaf_83_clk),
    .Q(\u0.subword[15] ),
    .QN(_00424_));
 DFF_X1 \u0.u3.d[0]$_DFF_P_  (.D(_00024_),
    .CK(clknet_leaf_28_clk),
    .Q(\u0.subword[0] ),
    .QN(_00411_));
 DFF_X1 \u0.u3.d[1]$_DFF_P_  (.D(_00025_),
    .CK(clknet_leaf_24_clk),
    .Q(\u0.subword[1] ),
    .QN(_00412_));
 DFF_X1 \u0.u3.d[2]$_DFF_P_  (.D(_00026_),
    .CK(clknet_leaf_23_clk),
    .Q(\u0.subword[2] ),
    .QN(_00409_));
 DFF_X1 \u0.u3.d[3]$_DFF_P_  (.D(_00027_),
    .CK(clknet_leaf_23_clk),
    .Q(\u0.subword[3] ),
    .QN(_00413_));
 DFF_X1 \u0.u3.d[4]$_DFF_P_  (.D(_00028_),
    .CK(clknet_leaf_35_clk),
    .Q(\u0.subword[4] ),
    .QN(_00414_));
 DFF_X1 \u0.u3.d[5]$_DFF_P_  (.D(_00029_),
    .CK(clknet_leaf_33_clk),
    .Q(\u0.subword[5] ),
    .QN(_00415_));
 DFF_X1 \u0.u3.d[6]$_DFF_P_  (.D(_00030_),
    .CK(clknet_leaf_36_clk),
    .Q(\u0.subword[6] ),
    .QN(_00416_));
 DFF_X1 \u0.u3.d[7]$_DFF_P_  (.D(_00031_),
    .CK(clknet_leaf_32_clk),
    .Q(\u0.subword[7] ),
    .QN(_00417_));
 DFF_X1 \u0.w[0][0]$_DFF_P_  (.D(_00289_),
    .CK(clknet_leaf_31_clk),
    .Q(\u0.w[0][0] ),
    .QN(_14531_));
 DFF_X1 \u0.w[0][10]$_DFF_P_  (.D(_00290_),
    .CK(clknet_leaf_24_clk),
    .Q(\u0.w[0][10] ),
    .QN(_14532_));
 DFF_X1 \u0.w[0][11]$_DFF_P_  (.D(_00291_),
    .CK(clknet_leaf_80_clk),
    .Q(\u0.w[0][11] ),
    .QN(_14533_));
 DFF_X1 \u0.w[0][12]$_DFF_P_  (.D(_00292_),
    .CK(clknet_leaf_78_clk),
    .Q(\u0.w[0][12] ),
    .QN(_14534_));
 DFF_X1 \u0.w[0][13]$_DFF_P_  (.D(_00293_),
    .CK(clknet_leaf_80_clk),
    .Q(\u0.w[0][13] ),
    .QN(_14535_));
 DFF_X1 \u0.w[0][14]$_DFF_P_  (.D(_00294_),
    .CK(clknet_leaf_7_clk),
    .Q(\u0.w[0][14] ),
    .QN(_14536_));
 DFF_X1 \u0.w[0][15]$_DFF_P_  (.D(_00295_),
    .CK(clknet_leaf_76_clk),
    .Q(\u0.w[0][15] ),
    .QN(_14537_));
 DFF_X1 \u0.w[0][16]$_DFF_P_  (.D(_00296_),
    .CK(clknet_leaf_6_clk),
    .Q(\u0.w[0][16] ),
    .QN(_14538_));
 DFF_X1 \u0.w[0][17]$_DFF_P_  (.D(_00297_),
    .CK(clknet_leaf_86_clk),
    .Q(\u0.w[0][17] ),
    .QN(_14539_));
 DFF_X1 \u0.w[0][18]$_DFF_P_  (.D(_00298_),
    .CK(clknet_leaf_81_clk),
    .Q(\u0.w[0][18] ),
    .QN(_14540_));
 DFF_X1 \u0.w[0][19]$_DFF_P_  (.D(_00299_),
    .CK(clknet_leaf_81_clk),
    .Q(\u0.w[0][19] ),
    .QN(_14541_));
 DFF_X1 \u0.w[0][1]$_DFF_P_  (.D(_00300_),
    .CK(clknet_leaf_37_clk),
    .Q(\u0.w[0][1] ),
    .QN(_14542_));
 DFF_X1 \u0.w[0][20]$_DFF_P_  (.D(_00301_),
    .CK(clknet_leaf_90_clk),
    .Q(\u0.w[0][20] ),
    .QN(_14543_));
 DFF_X1 \u0.w[0][21]$_DFF_P_  (.D(_00302_),
    .CK(clknet_leaf_84_clk),
    .Q(\u0.w[0][21] ),
    .QN(_14544_));
 DFF_X1 \u0.w[0][22]$_DFF_P_  (.D(_00303_),
    .CK(clknet_leaf_85_clk),
    .Q(\u0.w[0][22] ),
    .QN(_14545_));
 DFF_X1 \u0.w[0][23]$_DFF_P_  (.D(_00304_),
    .CK(clknet_leaf_84_clk),
    .Q(\u0.w[0][23] ),
    .QN(_14546_));
 DFF_X1 \u0.w[0][24]$_DFF_P_  (.D(_00305_),
    .CK(clknet_leaf_80_clk),
    .Q(\u0.w[0][24] ),
    .QN(_14547_));
 DFF_X1 \u0.w[0][25]$_DFF_P_  (.D(_00306_),
    .CK(clknet_leaf_79_clk),
    .Q(\u0.w[0][25] ),
    .QN(_14548_));
 DFF_X1 \u0.w[0][26]$_DFF_P_  (.D(_00307_),
    .CK(clknet_leaf_78_clk),
    .Q(\u0.w[0][26] ),
    .QN(_14549_));
 DFF_X1 \u0.w[0][27]$_DFF_P_  (.D(_00308_),
    .CK(clknet_leaf_78_clk),
    .Q(\u0.w[0][27] ),
    .QN(_14550_));
 DFF_X1 \u0.w[0][28]$_DFF_P_  (.D(_00309_),
    .CK(clknet_leaf_83_clk),
    .Q(\u0.w[0][28] ),
    .QN(_14551_));
 DFF_X1 \u0.w[0][29]$_DFF_P_  (.D(_00310_),
    .CK(clknet_leaf_83_clk),
    .Q(\u0.w[0][29] ),
    .QN(_14552_));
 DFF_X1 \u0.w[0][2]$_DFF_P_  (.D(_00311_),
    .CK(clknet_leaf_23_clk),
    .Q(\u0.w[0][2] ),
    .QN(_14553_));
 DFF_X1 \u0.w[0][30]$_DFF_P_  (.D(_00312_),
    .CK(clknet_leaf_83_clk),
    .Q(\u0.w[0][30] ),
    .QN(_14554_));
 DFF_X1 \u0.w[0][31]$_DFF_P_  (.D(_00313_),
    .CK(clknet_leaf_76_clk),
    .Q(\u0.w[0][31] ),
    .QN(_14555_));
 DFF_X1 \u0.w[0][3]$_DFF_P_  (.D(_00314_),
    .CK(clknet_leaf_37_clk),
    .Q(\u0.w[0][3] ),
    .QN(_14556_));
 DFF_X1 \u0.w[0][4]$_DFF_P_  (.D(_00315_),
    .CK(clknet_leaf_34_clk),
    .Q(\u0.w[0][4] ),
    .QN(_14557_));
 DFF_X1 \u0.w[0][5]$_DFF_P_  (.D(_00316_),
    .CK(clknet_leaf_51_clk),
    .Q(\u0.w[0][5] ),
    .QN(_14558_));
 DFF_X1 \u0.w[0][6]$_DFF_P_  (.D(_00317_),
    .CK(clknet_leaf_35_clk),
    .Q(\u0.w[0][6] ),
    .QN(_14559_));
 DFF_X1 \u0.w[0][7]$_DFF_P_  (.D(_00318_),
    .CK(clknet_leaf_31_clk),
    .Q(\u0.w[0][7] ),
    .QN(_14560_));
 DFF_X1 \u0.w[0][8]$_DFF_P_  (.D(_00319_),
    .CK(clknet_leaf_27_clk),
    .Q(\u0.w[0][8] ),
    .QN(_14561_));
 DFF_X1 \u0.w[0][9]$_DFF_P_  (.D(_00320_),
    .CK(clknet_leaf_27_clk),
    .Q(\u0.w[0][9] ),
    .QN(_14562_));
 DFF_X1 \u0.w[1][0]$_DFF_P_  (.D(_00321_),
    .CK(clknet_leaf_31_clk),
    .Q(\u0.w[1][0] ),
    .QN(_14563_));
 DFF_X1 \u0.w[1][10]$_DFF_P_  (.D(_00322_),
    .CK(clknet_leaf_77_clk),
    .Q(\u0.w[1][10] ),
    .QN(_14564_));
 DFF_X1 \u0.w[1][11]$_DFF_P_  (.D(_00323_),
    .CK(clknet_leaf_78_clk),
    .Q(\u0.w[1][11] ),
    .QN(_14565_));
 DFF_X1 \u0.w[1][12]$_DFF_P_  (.D(_00324_),
    .CK(clknet_leaf_78_clk),
    .Q(\u0.w[1][12] ),
    .QN(_14566_));
 DFF_X1 \u0.w[1][13]$_DFF_P_  (.D(_00325_),
    .CK(clknet_leaf_79_clk),
    .Q(\u0.w[1][13] ),
    .QN(_14567_));
 DFF_X1 \u0.w[1][14]$_DFF_P_  (.D(_00326_),
    .CK(clknet_leaf_7_clk),
    .Q(\u0.w[1][14] ),
    .QN(_14568_));
 DFF_X1 \u0.w[1][15]$_DFF_P_  (.D(_00327_),
    .CK(clknet_leaf_83_clk),
    .Q(\u0.w[1][15] ),
    .QN(_14569_));
 DFF_X1 \u0.w[1][16]$_DFF_P_  (.D(_00328_),
    .CK(clknet_leaf_6_clk),
    .Q(\u0.w[1][16] ),
    .QN(_14570_));
 DFF_X1 \u0.w[1][17]$_DFF_P_  (.D(_00329_),
    .CK(clknet_leaf_81_clk),
    .Q(\u0.w[1][17] ),
    .QN(_14571_));
 DFF_X1 \u0.w[1][18]$_DFF_P_  (.D(_00330_),
    .CK(clknet_leaf_80_clk),
    .Q(\u0.w[1][18] ),
    .QN(_14572_));
 DFF_X1 \u0.w[1][19]$_DFF_P_  (.D(_00331_),
    .CK(clknet_leaf_81_clk),
    .Q(\u0.w[1][19] ),
    .QN(_14573_));
 DFF_X1 \u0.w[1][1]$_DFF_P_  (.D(_00332_),
    .CK(clknet_leaf_37_clk),
    .Q(\u0.w[1][1] ),
    .QN(_14574_));
 DFF_X1 \u0.w[1][20]$_DFF_P_  (.D(_00333_),
    .CK(clknet_leaf_85_clk),
    .Q(\u0.w[1][20] ),
    .QN(_14575_));
 DFF_X1 \u0.w[1][21]$_DFF_P_  (.D(_00334_),
    .CK(clknet_leaf_84_clk),
    .Q(\u0.w[1][21] ),
    .QN(_14576_));
 DFF_X1 \u0.w[1][22]$_DFF_P_  (.D(_00335_),
    .CK(clknet_leaf_86_clk),
    .Q(\u0.w[1][22] ),
    .QN(_14577_));
 DFF_X1 \u0.w[1][23]$_DFF_P_  (.D(_00336_),
    .CK(clknet_leaf_82_clk),
    .Q(\u0.w[1][23] ),
    .QN(_14578_));
 DFF_X1 \u0.w[1][24]$_DFF_P_  (.D(_00337_),
    .CK(clknet_leaf_53_clk),
    .Q(\u0.w[1][24] ),
    .QN(_14579_));
 DFF_X1 \u0.w[1][25]$_DFF_P_  (.D(_00338_),
    .CK(clknet_leaf_47_clk),
    .Q(\u0.w[1][25] ),
    .QN(_14580_));
 DFF_X1 \u0.w[1][26]$_DFF_P_  (.D(_00339_),
    .CK(clknet_leaf_57_clk),
    .Q(\u0.w[1][26] ),
    .QN(_14581_));
 DFF_X1 \u0.w[1][27]$_DFF_P_  (.D(_00340_),
    .CK(clknet_leaf_62_clk),
    .Q(\u0.w[1][27] ),
    .QN(_14582_));
 DFF_X1 \u0.w[1][28]$_DFF_P_  (.D(_00341_),
    .CK(clknet_leaf_63_clk),
    .Q(\u0.w[1][28] ),
    .QN(_14583_));
 DFF_X1 \u0.w[1][29]$_DFF_P_  (.D(_00342_),
    .CK(clknet_leaf_63_clk),
    .Q(\u0.w[1][29] ),
    .QN(_14584_));
 DFF_X1 \u0.w[1][2]$_DFF_P_  (.D(_00343_),
    .CK(clknet_leaf_23_clk),
    .Q(\u0.w[1][2] ),
    .QN(_14585_));
 DFF_X1 \u0.w[1][30]$_DFF_P_  (.D(_00344_),
    .CK(clknet_leaf_63_clk),
    .Q(\u0.w[1][30] ),
    .QN(_14586_));
 DFF_X1 \u0.w[1][31]$_DFF_P_  (.D(_00345_),
    .CK(clknet_leaf_46_clk),
    .Q(\u0.w[1][31] ),
    .QN(_14587_));
 DFF_X1 \u0.w[1][3]$_DFF_P_  (.D(_00346_),
    .CK(clknet_leaf_36_clk),
    .Q(\u0.w[1][3] ),
    .QN(_14588_));
 DFF_X1 \u0.w[1][4]$_DFF_P_  (.D(_00347_),
    .CK(clknet_leaf_35_clk),
    .Q(\u0.w[1][4] ),
    .QN(_14589_));
 DFF_X1 \u0.w[1][5]$_DFF_P_  (.D(_00348_),
    .CK(clknet_leaf_33_clk),
    .Q(\u0.w[1][5] ),
    .QN(_14590_));
 DFF_X1 \u0.w[1][6]$_DFF_P_  (.D(_00349_),
    .CK(clknet_leaf_35_clk),
    .Q(\u0.w[1][6] ),
    .QN(_14591_));
 DFF_X1 \u0.w[1][7]$_DFF_P_  (.D(_00350_),
    .CK(clknet_leaf_32_clk),
    .Q(\u0.w[1][7] ),
    .QN(_14592_));
 DFF_X1 \u0.w[1][8]$_DFF_P_  (.D(_00351_),
    .CK(clknet_leaf_8_clk),
    .Q(\u0.w[1][8] ),
    .QN(_14593_));
 DFF_X1 \u0.w[1][9]$_DFF_P_  (.D(_00352_),
    .CK(clknet_leaf_8_clk),
    .Q(\u0.w[1][9] ),
    .QN(_14594_));
 DFF_X1 \u0.w[2][0]$_DFF_P_  (.D(_00353_),
    .CK(clknet_leaf_36_clk),
    .Q(\u0.w[2][0] ),
    .QN(_14595_));
 DFF_X1 \u0.w[2][10]$_DFF_P_  (.D(_00354_),
    .CK(clknet_leaf_77_clk),
    .Q(\u0.w[2][10] ),
    .QN(_14596_));
 DFF_X1 \u0.w[2][11]$_DFF_P_  (.D(_00355_),
    .CK(clknet_leaf_80_clk),
    .Q(\u0.w[2][11] ),
    .QN(_14597_));
 DFF_X1 \u0.w[2][12]$_DFF_P_  (.D(_00356_),
    .CK(clknet_leaf_79_clk),
    .Q(\u0.w[2][12] ),
    .QN(_14598_));
 DFF_X1 \u0.w[2][13]$_DFF_P_  (.D(_00357_),
    .CK(clknet_leaf_79_clk),
    .Q(\u0.w[2][13] ),
    .QN(_14599_));
 DFF_X1 \u0.w[2][14]$_DFF_P_  (.D(_00358_),
    .CK(clknet_leaf_78_clk),
    .Q(\u0.w[2][14] ),
    .QN(_14600_));
 DFF_X1 \u0.w[2][15]$_DFF_P_  (.D(_00359_),
    .CK(clknet_leaf_83_clk),
    .Q(\u0.w[2][15] ),
    .QN(_14601_));
 DFF_X1 \u0.w[2][16]$_DFF_P_  (.D(_00360_),
    .CK(clknet_leaf_80_clk),
    .Q(\u0.w[2][16] ),
    .QN(_14602_));
 DFF_X1 \u0.w[2][17]$_DFF_P_  (.D(_00361_),
    .CK(clknet_leaf_82_clk),
    .Q(\u0.w[2][17] ),
    .QN(_14603_));
 DFF_X1 \u0.w[2][18]$_DFF_P_  (.D(_00362_),
    .CK(clknet_leaf_6_clk),
    .Q(\u0.w[2][18] ),
    .QN(_14604_));
 DFF_X1 \u0.w[2][19]$_DFF_P_  (.D(_00363_),
    .CK(clknet_leaf_82_clk),
    .Q(\u0.w[2][19] ),
    .QN(_14605_));
 DFF_X1 \u0.w[2][1]$_DFF_P_  (.D(_00364_),
    .CK(clknet_leaf_36_clk),
    .Q(\u0.w[2][1] ),
    .QN(_14606_));
 DFF_X1 \u0.w[2][20]$_DFF_P_  (.D(_00365_),
    .CK(clknet_leaf_85_clk),
    .Q(\u0.w[2][20] ),
    .QN(_14607_));
 DFF_X1 \u0.w[2][21]$_DFF_P_  (.D(_00366_),
    .CK(clknet_leaf_91_clk),
    .Q(\u0.w[2][21] ),
    .QN(_14608_));
 DFF_X1 \u0.w[2][22]$_DFF_P_  (.D(_00367_),
    .CK(clknet_leaf_86_clk),
    .Q(\u0.w[2][22] ),
    .QN(_14609_));
 DFF_X1 \u0.w[2][23]$_DFF_P_  (.D(_00368_),
    .CK(clknet_leaf_82_clk),
    .Q(\u0.w[2][23] ),
    .QN(_14610_));
 DFF_X1 \u0.w[2][24]$_DFF_P_  (.D(_00369_),
    .CK(clknet_leaf_47_clk),
    .Q(\u0.w[2][24] ),
    .QN(_14611_));
 DFF_X1 \u0.w[2][25]$_DFF_P_  (.D(_00370_),
    .CK(clknet_leaf_47_clk),
    .Q(\u0.w[2][25] ),
    .QN(_14612_));
 DFF_X1 \u0.w[2][26]$_DFF_P_  (.D(_00371_),
    .CK(clknet_leaf_57_clk),
    .Q(\u0.w[2][26] ),
    .QN(_14613_));
 DFF_X1 \u0.w[2][27]$_DFF_P_  (.D(_00372_),
    .CK(clknet_leaf_63_clk),
    .Q(\u0.w[2][27] ),
    .QN(_14614_));
 DFF_X1 \u0.w[2][28]$_DFF_P_  (.D(_00373_),
    .CK(clknet_leaf_62_clk),
    .Q(\u0.w[2][28] ),
    .QN(_14615_));
 DFF_X1 \u0.w[2][29]$_DFF_P_  (.D(_00374_),
    .CK(clknet_leaf_63_clk),
    .Q(\u0.w[2][29] ),
    .QN(_14616_));
 DFF_X1 \u0.w[2][2]$_DFF_P_  (.D(_00375_),
    .CK(clknet_leaf_23_clk),
    .Q(\u0.w[2][2] ),
    .QN(_14617_));
 DFF_X1 \u0.w[2][30]$_DFF_P_  (.D(_00376_),
    .CK(clknet_leaf_63_clk),
    .Q(\u0.w[2][30] ),
    .QN(_14618_));
 DFF_X1 \u0.w[2][31]$_DFF_P_  (.D(_00377_),
    .CK(clknet_leaf_46_clk),
    .Q(\u0.w[2][31] ),
    .QN(_14619_));
 DFF_X1 \u0.w[2][3]$_DFF_P_  (.D(_00378_),
    .CK(clknet_leaf_36_clk),
    .Q(\u0.w[2][3] ),
    .QN(_14620_));
 DFF_X1 \u0.w[2][4]$_DFF_P_  (.D(_00379_),
    .CK(clknet_leaf_34_clk),
    .Q(\u0.w[2][4] ),
    .QN(_14621_));
 DFF_X1 \u0.w[2][5]$_DFF_P_  (.D(_00380_),
    .CK(clknet_leaf_51_clk),
    .Q(\u0.w[2][5] ),
    .QN(_14622_));
 DFF_X1 \u0.w[2][6]$_DFF_P_  (.D(_00381_),
    .CK(clknet_leaf_35_clk),
    .Q(\u0.w[2][6] ),
    .QN(_14623_));
 DFF_X1 \u0.w[2][7]$_DFF_P_  (.D(_00382_),
    .CK(clknet_leaf_32_clk),
    .Q(\u0.w[2][7] ),
    .QN(_14624_));
 DFF_X1 \u0.w[2][8]$_DFF_P_  (.D(_00383_),
    .CK(clknet_leaf_8_clk),
    .Q(\u0.w[2][8] ),
    .QN(_14625_));
 DFF_X1 \u0.w[2][9]$_DFF_P_  (.D(_00384_),
    .CK(clknet_leaf_8_clk),
    .Q(\u0.w[2][9] ),
    .QN(_14626_));
 DFF_X1 \u0.w[3][0]$_DFF_P_  (.D(net49),
    .CK(clknet_leaf_24_clk),
    .Q(\u0.tmp_w[0] ),
    .QN(_14627_));
 DFF_X1 \u0.w[3][10]$_DFF_P_  (.D(_14717_),
    .CK(clknet_leaf_2_clk),
    .Q(\u0.tmp_w[10] ),
    .QN(_14628_));
 DFF_X1 \u0.w[3][11]$_DFF_P_  (.D(_00385_),
    .CK(clknet_leaf_2_clk),
    .Q(\u0.tmp_w[11] ),
    .QN(_14629_));
 DFF_X1 \u0.w[3][12]$_DFF_P_  (.D(_00386_),
    .CK(clknet_leaf_2_clk),
    .Q(\u0.tmp_w[12] ),
    .QN(_14630_));
 DFF_X1 \u0.w[3][13]$_DFF_P_  (.D(_00387_),
    .CK(clknet_leaf_2_clk),
    .Q(\u0.tmp_w[13] ),
    .QN(_14631_));
 DFF_X1 \u0.w[3][14]$_DFF_P_  (.D(_00388_),
    .CK(clknet_leaf_1_clk),
    .Q(\u0.tmp_w[14] ),
    .QN(_14632_));
 DFF_X1 \u0.w[3][15]$_DFF_P_  (.D(_00389_),
    .CK(clknet_leaf_3_clk),
    .Q(\u0.tmp_w[15] ),
    .QN(_14633_));
 DFF_X1 \u0.w[3][16]$_DFF_P_  (.D(net801),
    .CK(clknet_leaf_88_clk),
    .Q(\u0.tmp_w[16] ),
    .QN(_14634_));
 DFF_X1 \u0.w[3][17]$_DFF_P_  (.D(net66),
    .CK(clknet_leaf_95_clk),
    .Q(\u0.tmp_w[17] ),
    .QN(_14635_));
 DFF_X1 \u0.w[3][18]$_DFF_P_  (.D(_14683_),
    .CK(clknet_leaf_90_clk),
    .Q(\u0.tmp_w[18] ),
    .QN(_14636_));
 DFF_X1 \u0.w[3][19]$_DFF_P_  (.D(_00390_),
    .CK(clknet_leaf_89_clk),
    .Q(\u0.tmp_w[19] ),
    .QN(_14637_));
 DFF_X1 \u0.w[3][1]$_DFF_P_  (.D(net27),
    .CK(clknet_leaf_25_clk),
    .Q(\u0.tmp_w[1] ),
    .QN(_14638_));
 DFF_X1 \u0.w[3][20]$_DFF_P_  (.D(_00391_),
    .CK(clknet_leaf_89_clk),
    .Q(\u0.tmp_w[20] ),
    .QN(_14639_));
 DFF_X1 \u0.w[3][21]$_DFF_P_  (.D(_00392_),
    .CK(clknet_leaf_89_clk),
    .Q(\u0.tmp_w[21] ),
    .QN(_14640_));
 DFF_X1 \u0.w[3][22]$_DFF_P_  (.D(_00393_),
    .CK(clknet_leaf_95_clk),
    .Q(\u0.tmp_w[22] ),
    .QN(_14641_));
 DFF_X1 \u0.w[3][23]$_DFF_P_  (.D(_00394_),
    .CK(clknet_leaf_88_clk),
    .Q(\u0.tmp_w[23] ),
    .QN(_14642_));
 DFF_X1 \u0.w[3][24]$_DFF_P_  (.D(_14761_),
    .CK(clknet_leaf_15_clk),
    .Q(\u0.tmp_w[24] ),
    .QN(_14643_));
 DFF_X1 \u0.w[3][25]$_DFF_P_  (.D(_14760_),
    .CK(clknet_leaf_16_clk),
    .Q(\u0.tmp_w[25] ),
    .QN(_14644_));
 DFF_X1 \u0.w[3][26]$_DFF_P_  (.D(_14780_),
    .CK(clknet_leaf_14_clk),
    .Q(\u0.tmp_w[26] ),
    .QN(_14645_));
 DFF_X1 \u0.w[3][27]$_DFF_P_  (.D(_00395_),
    .CK(clknet_leaf_14_clk),
    .Q(\u0.tmp_w[27] ),
    .QN(_14646_));
 DFF_X1 \u0.w[3][28]$_DFF_P_  (.D(_00396_),
    .CK(clknet_leaf_27_clk),
    .Q(\u0.tmp_w[28] ),
    .QN(_14647_));
 DFF_X1 \u0.w[3][29]$_DFF_P_  (.D(_00397_),
    .CK(clknet_leaf_15_clk),
    .Q(\u0.tmp_w[29] ),
    .QN(_14648_));
 DFF_X1 \u0.w[3][2]$_DFF_P_  (.D(_14751_),
    .CK(clknet_leaf_24_clk),
    .Q(\u0.tmp_w[2] ),
    .QN(_14649_));
 DFF_X1 \u0.w[3][30]$_DFF_P_  (.D(_00398_),
    .CK(clknet_leaf_11_clk),
    .Q(\u0.tmp_w[30] ),
    .QN(_14650_));
 DFF_X1 \u0.w[3][31]$_DFF_P_  (.D(_00399_),
    .CK(clknet_leaf_15_clk),
    .Q(\u0.tmp_w[31] ),
    .QN(_14651_));
 DFF_X1 \u0.w[3][3]$_DFF_P_  (.D(_00400_),
    .CK(clknet_leaf_26_clk),
    .Q(\u0.tmp_w[3] ),
    .QN(_14652_));
 DFF_X1 \u0.w[3][4]$_DFF_P_  (.D(_00401_),
    .CK(clknet_leaf_26_clk),
    .Q(\u0.tmp_w[4] ),
    .QN(_14653_));
 DFF_X1 \u0.w[3][5]$_DFF_P_  (.D(_00402_),
    .CK(clknet_leaf_25_clk),
    .Q(\u0.tmp_w[5] ),
    .QN(_14654_));
 DFF_X1 \u0.w[3][6]$_DFF_P_  (.D(_00403_),
    .CK(clknet_leaf_25_clk),
    .Q(\u0.tmp_w[6] ),
    .QN(_14655_));
 DFF_X2 \u0.w[3][7]$_DFF_P_  (.D(_00404_),
    .CK(clknet_leaf_25_clk),
    .Q(\u0.tmp_w[7] ),
    .QN(_14656_));
 DFF_X1 \u0.w[3][8]$_DFF_P_  (.D(_14693_),
    .CK(clknet_leaf_2_clk),
    .Q(\u0.tmp_w[8] ),
    .QN(_14657_));
 DFF_X1 \u0.w[3][9]$_DFF_P_  (.D(net14),
    .CK(clknet_leaf_1_clk),
    .Q(\u0.tmp_w[9] ),
    .QN(_14178_));
 BUF_X4 clone103 (.A(_05531_),
    .Z(net103));
 BUF_X8 clone105 (.A(_05709_),
    .Z(net105));
 BUF_X8 split111 (.A(net485),
    .Z(net111));
 BUF_X4 clone112 (.A(_09734_),
    .Z(net112));
 BUF_X4 clone113 (.A(_09735_),
    .Z(net113));
 BUF_X8 clone114 (.A(_09736_),
    .Z(net114));
 INV_X2 clone123 (.A(net124),
    .ZN(net123));
 NOR2_X4 clone124 (.A1(_09001_),
    .A2(_08991_),
    .ZN(net124));
 NOR2_X4 clone125 (.A1(_01602_),
    .A2(net592),
    .ZN(net125));
 BUF_X2 clone175 (.A(_15002_),
    .Z(net175));
 BUF_X4 clone176 (.A(_13176_),
    .Z(net176));
 BUF_X4 clone177 (.A(_13177_),
    .Z(net177));
 BUF_X8 clone178 (.A(_13178_),
    .Z(net178));
 TAPCELL_X1 PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Right_29 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Right_30 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Right_31 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Right_32 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Right_33 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Right_34 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Right_35 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Right_36 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Right_37 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Right_38 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Right_39 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Right_40 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Right_41 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Right_42 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Right_43 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Right_44 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Right_45 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Right_46 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Right_47 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Right_48 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Right_49 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Right_50 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Right_51 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Right_52 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Right_53 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Right_54 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Right_55 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Right_56 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Right_57 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Right_58 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Right_59 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Right_60 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Right_61 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Right_62 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Right_63 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Right_64 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Right_65 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Right_66 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Right_67 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Right_68 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Right_69 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Right_70 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Right_71 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Right_72 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Right_73 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Right_74 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Right_75 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Right_76 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Right_77 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Right_78 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Right_79 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Right_80 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Right_81 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Right_82 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Right_83 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Right_84 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Right_85 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Right_86 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Right_87 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Right_88 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Right_89 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Right_90 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Right_91 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Right_92 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Right_93 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Right_94 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Right_95 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Right_96 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Right_97 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Right_98 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Right_99 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Right_100 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Right_101 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Right_102 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Right_103 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Right_104 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Right_105 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Right_106 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Right_107 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Right_108 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Right_109 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Right_110 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Right_111 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Right_112 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Right_113 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Right_114 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Right_115 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Right_116 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Right_117 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Right_118 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Right_119 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Right_120 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Right_121 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Right_122 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Right_123 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Right_124 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Right_125 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Right_126 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Right_127 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Right_128 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Right_129 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Right_130 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Right_131 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Right_132 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Right_133 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Right_134 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Right_135 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Right_136 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Right_137 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Right_138 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Right_139 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Right_140 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Right_141 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Right_142 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Right_143 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Right_144 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Right_145 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Right_146 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Right_147 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Right_148 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Right_149 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Right_150 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Right_151 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Right_152 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Right_153 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Right_154 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Right_155 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Right_156 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Right_157 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Right_158 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Right_159 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Right_160 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Right_161 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Right_162 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Right_163 ();
 TAPCELL_X1 PHY_EDGE_ROW_0_Left_164 ();
 TAPCELL_X1 PHY_EDGE_ROW_1_Left_165 ();
 TAPCELL_X1 PHY_EDGE_ROW_2_Left_166 ();
 TAPCELL_X1 PHY_EDGE_ROW_3_Left_167 ();
 TAPCELL_X1 PHY_EDGE_ROW_4_Left_168 ();
 TAPCELL_X1 PHY_EDGE_ROW_5_Left_169 ();
 TAPCELL_X1 PHY_EDGE_ROW_6_Left_170 ();
 TAPCELL_X1 PHY_EDGE_ROW_7_Left_171 ();
 TAPCELL_X1 PHY_EDGE_ROW_8_Left_172 ();
 TAPCELL_X1 PHY_EDGE_ROW_9_Left_173 ();
 TAPCELL_X1 PHY_EDGE_ROW_10_Left_174 ();
 TAPCELL_X1 PHY_EDGE_ROW_11_Left_175 ();
 TAPCELL_X1 PHY_EDGE_ROW_12_Left_176 ();
 TAPCELL_X1 PHY_EDGE_ROW_13_Left_177 ();
 TAPCELL_X1 PHY_EDGE_ROW_14_Left_178 ();
 TAPCELL_X1 PHY_EDGE_ROW_15_Left_179 ();
 TAPCELL_X1 PHY_EDGE_ROW_16_Left_180 ();
 TAPCELL_X1 PHY_EDGE_ROW_17_Left_181 ();
 TAPCELL_X1 PHY_EDGE_ROW_18_Left_182 ();
 TAPCELL_X1 PHY_EDGE_ROW_19_Left_183 ();
 TAPCELL_X1 PHY_EDGE_ROW_20_Left_184 ();
 TAPCELL_X1 PHY_EDGE_ROW_21_Left_185 ();
 TAPCELL_X1 PHY_EDGE_ROW_22_Left_186 ();
 TAPCELL_X1 PHY_EDGE_ROW_23_Left_187 ();
 TAPCELL_X1 PHY_EDGE_ROW_24_Left_188 ();
 TAPCELL_X1 PHY_EDGE_ROW_25_Left_189 ();
 TAPCELL_X1 PHY_EDGE_ROW_26_Left_190 ();
 TAPCELL_X1 PHY_EDGE_ROW_27_Left_191 ();
 TAPCELL_X1 PHY_EDGE_ROW_28_Left_192 ();
 TAPCELL_X1 PHY_EDGE_ROW_29_Left_193 ();
 TAPCELL_X1 PHY_EDGE_ROW_30_Left_194 ();
 TAPCELL_X1 PHY_EDGE_ROW_31_Left_195 ();
 TAPCELL_X1 PHY_EDGE_ROW_32_Left_196 ();
 TAPCELL_X1 PHY_EDGE_ROW_33_Left_197 ();
 TAPCELL_X1 PHY_EDGE_ROW_34_Left_198 ();
 TAPCELL_X1 PHY_EDGE_ROW_35_Left_199 ();
 TAPCELL_X1 PHY_EDGE_ROW_36_Left_200 ();
 TAPCELL_X1 PHY_EDGE_ROW_37_Left_201 ();
 TAPCELL_X1 PHY_EDGE_ROW_38_Left_202 ();
 TAPCELL_X1 PHY_EDGE_ROW_39_Left_203 ();
 TAPCELL_X1 PHY_EDGE_ROW_40_Left_204 ();
 TAPCELL_X1 PHY_EDGE_ROW_41_Left_205 ();
 TAPCELL_X1 PHY_EDGE_ROW_42_Left_206 ();
 TAPCELL_X1 PHY_EDGE_ROW_43_Left_207 ();
 TAPCELL_X1 PHY_EDGE_ROW_44_Left_208 ();
 TAPCELL_X1 PHY_EDGE_ROW_45_Left_209 ();
 TAPCELL_X1 PHY_EDGE_ROW_46_Left_210 ();
 TAPCELL_X1 PHY_EDGE_ROW_47_Left_211 ();
 TAPCELL_X1 PHY_EDGE_ROW_48_Left_212 ();
 TAPCELL_X1 PHY_EDGE_ROW_49_Left_213 ();
 TAPCELL_X1 PHY_EDGE_ROW_50_Left_214 ();
 TAPCELL_X1 PHY_EDGE_ROW_51_Left_215 ();
 TAPCELL_X1 PHY_EDGE_ROW_52_Left_216 ();
 TAPCELL_X1 PHY_EDGE_ROW_53_Left_217 ();
 TAPCELL_X1 PHY_EDGE_ROW_54_Left_218 ();
 TAPCELL_X1 PHY_EDGE_ROW_55_Left_219 ();
 TAPCELL_X1 PHY_EDGE_ROW_56_Left_220 ();
 TAPCELL_X1 PHY_EDGE_ROW_57_Left_221 ();
 TAPCELL_X1 PHY_EDGE_ROW_58_Left_222 ();
 TAPCELL_X1 PHY_EDGE_ROW_59_Left_223 ();
 TAPCELL_X1 PHY_EDGE_ROW_60_Left_224 ();
 TAPCELL_X1 PHY_EDGE_ROW_61_Left_225 ();
 TAPCELL_X1 PHY_EDGE_ROW_62_Left_226 ();
 TAPCELL_X1 PHY_EDGE_ROW_63_Left_227 ();
 TAPCELL_X1 PHY_EDGE_ROW_64_Left_228 ();
 TAPCELL_X1 PHY_EDGE_ROW_65_Left_229 ();
 TAPCELL_X1 PHY_EDGE_ROW_66_Left_230 ();
 TAPCELL_X1 PHY_EDGE_ROW_67_Left_231 ();
 TAPCELL_X1 PHY_EDGE_ROW_68_Left_232 ();
 TAPCELL_X1 PHY_EDGE_ROW_69_Left_233 ();
 TAPCELL_X1 PHY_EDGE_ROW_70_Left_234 ();
 TAPCELL_X1 PHY_EDGE_ROW_71_Left_235 ();
 TAPCELL_X1 PHY_EDGE_ROW_72_Left_236 ();
 TAPCELL_X1 PHY_EDGE_ROW_73_Left_237 ();
 TAPCELL_X1 PHY_EDGE_ROW_74_Left_238 ();
 TAPCELL_X1 PHY_EDGE_ROW_75_Left_239 ();
 TAPCELL_X1 PHY_EDGE_ROW_76_Left_240 ();
 TAPCELL_X1 PHY_EDGE_ROW_77_Left_241 ();
 TAPCELL_X1 PHY_EDGE_ROW_78_Left_242 ();
 TAPCELL_X1 PHY_EDGE_ROW_79_Left_243 ();
 TAPCELL_X1 PHY_EDGE_ROW_80_Left_244 ();
 TAPCELL_X1 PHY_EDGE_ROW_81_Left_245 ();
 TAPCELL_X1 PHY_EDGE_ROW_82_Left_246 ();
 TAPCELL_X1 PHY_EDGE_ROW_83_Left_247 ();
 TAPCELL_X1 PHY_EDGE_ROW_84_Left_248 ();
 TAPCELL_X1 PHY_EDGE_ROW_85_Left_249 ();
 TAPCELL_X1 PHY_EDGE_ROW_86_Left_250 ();
 TAPCELL_X1 PHY_EDGE_ROW_87_Left_251 ();
 TAPCELL_X1 PHY_EDGE_ROW_88_Left_252 ();
 TAPCELL_X1 PHY_EDGE_ROW_89_Left_253 ();
 TAPCELL_X1 PHY_EDGE_ROW_90_Left_254 ();
 TAPCELL_X1 PHY_EDGE_ROW_91_Left_255 ();
 TAPCELL_X1 PHY_EDGE_ROW_92_Left_256 ();
 TAPCELL_X1 PHY_EDGE_ROW_93_Left_257 ();
 TAPCELL_X1 PHY_EDGE_ROW_94_Left_258 ();
 TAPCELL_X1 PHY_EDGE_ROW_95_Left_259 ();
 TAPCELL_X1 PHY_EDGE_ROW_96_Left_260 ();
 TAPCELL_X1 PHY_EDGE_ROW_97_Left_261 ();
 TAPCELL_X1 PHY_EDGE_ROW_98_Left_262 ();
 TAPCELL_X1 PHY_EDGE_ROW_99_Left_263 ();
 TAPCELL_X1 PHY_EDGE_ROW_100_Left_264 ();
 TAPCELL_X1 PHY_EDGE_ROW_101_Left_265 ();
 TAPCELL_X1 PHY_EDGE_ROW_102_Left_266 ();
 TAPCELL_X1 PHY_EDGE_ROW_103_Left_267 ();
 TAPCELL_X1 PHY_EDGE_ROW_104_Left_268 ();
 TAPCELL_X1 PHY_EDGE_ROW_105_Left_269 ();
 TAPCELL_X1 PHY_EDGE_ROW_106_Left_270 ();
 TAPCELL_X1 PHY_EDGE_ROW_107_Left_271 ();
 TAPCELL_X1 PHY_EDGE_ROW_108_Left_272 ();
 TAPCELL_X1 PHY_EDGE_ROW_109_Left_273 ();
 TAPCELL_X1 PHY_EDGE_ROW_110_Left_274 ();
 TAPCELL_X1 PHY_EDGE_ROW_111_Left_275 ();
 TAPCELL_X1 PHY_EDGE_ROW_112_Left_276 ();
 TAPCELL_X1 PHY_EDGE_ROW_113_Left_277 ();
 TAPCELL_X1 PHY_EDGE_ROW_114_Left_278 ();
 TAPCELL_X1 PHY_EDGE_ROW_115_Left_279 ();
 TAPCELL_X1 PHY_EDGE_ROW_116_Left_280 ();
 TAPCELL_X1 PHY_EDGE_ROW_117_Left_281 ();
 TAPCELL_X1 PHY_EDGE_ROW_118_Left_282 ();
 TAPCELL_X1 PHY_EDGE_ROW_119_Left_283 ();
 TAPCELL_X1 PHY_EDGE_ROW_120_Left_284 ();
 TAPCELL_X1 PHY_EDGE_ROW_121_Left_285 ();
 TAPCELL_X1 PHY_EDGE_ROW_122_Left_286 ();
 TAPCELL_X1 PHY_EDGE_ROW_123_Left_287 ();
 TAPCELL_X1 PHY_EDGE_ROW_124_Left_288 ();
 TAPCELL_X1 PHY_EDGE_ROW_125_Left_289 ();
 TAPCELL_X1 PHY_EDGE_ROW_126_Left_290 ();
 TAPCELL_X1 PHY_EDGE_ROW_127_Left_291 ();
 TAPCELL_X1 PHY_EDGE_ROW_128_Left_292 ();
 TAPCELL_X1 PHY_EDGE_ROW_129_Left_293 ();
 TAPCELL_X1 PHY_EDGE_ROW_130_Left_294 ();
 TAPCELL_X1 PHY_EDGE_ROW_131_Left_295 ();
 TAPCELL_X1 PHY_EDGE_ROW_132_Left_296 ();
 TAPCELL_X1 PHY_EDGE_ROW_133_Left_297 ();
 TAPCELL_X1 PHY_EDGE_ROW_134_Left_298 ();
 TAPCELL_X1 PHY_EDGE_ROW_135_Left_299 ();
 TAPCELL_X1 PHY_EDGE_ROW_136_Left_300 ();
 TAPCELL_X1 PHY_EDGE_ROW_137_Left_301 ();
 TAPCELL_X1 PHY_EDGE_ROW_138_Left_302 ();
 TAPCELL_X1 PHY_EDGE_ROW_139_Left_303 ();
 TAPCELL_X1 PHY_EDGE_ROW_140_Left_304 ();
 TAPCELL_X1 PHY_EDGE_ROW_141_Left_305 ();
 TAPCELL_X1 PHY_EDGE_ROW_142_Left_306 ();
 TAPCELL_X1 PHY_EDGE_ROW_143_Left_307 ();
 TAPCELL_X1 PHY_EDGE_ROW_144_Left_308 ();
 TAPCELL_X1 PHY_EDGE_ROW_145_Left_309 ();
 TAPCELL_X1 PHY_EDGE_ROW_146_Left_310 ();
 TAPCELL_X1 PHY_EDGE_ROW_147_Left_311 ();
 TAPCELL_X1 PHY_EDGE_ROW_148_Left_312 ();
 TAPCELL_X1 PHY_EDGE_ROW_149_Left_313 ();
 TAPCELL_X1 PHY_EDGE_ROW_150_Left_314 ();
 TAPCELL_X1 PHY_EDGE_ROW_151_Left_315 ();
 TAPCELL_X1 PHY_EDGE_ROW_152_Left_316 ();
 TAPCELL_X1 PHY_EDGE_ROW_153_Left_317 ();
 TAPCELL_X1 PHY_EDGE_ROW_154_Left_318 ();
 TAPCELL_X1 PHY_EDGE_ROW_155_Left_319 ();
 TAPCELL_X1 PHY_EDGE_ROW_156_Left_320 ();
 TAPCELL_X1 PHY_EDGE_ROW_157_Left_321 ();
 TAPCELL_X1 PHY_EDGE_ROW_158_Left_322 ();
 TAPCELL_X1 PHY_EDGE_ROW_159_Left_323 ();
 TAPCELL_X1 PHY_EDGE_ROW_160_Left_324 ();
 TAPCELL_X1 PHY_EDGE_ROW_161_Left_325 ();
 TAPCELL_X1 PHY_EDGE_ROW_162_Left_326 ();
 TAPCELL_X1 PHY_EDGE_ROW_163_Left_327 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_0_328 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_2_329 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_4_330 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_6_331 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_8_332 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_10_333 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_12_334 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_14_335 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_16_336 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_18_337 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_20_338 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_22_339 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_24_340 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_26_341 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_28_342 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_30_343 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_32_344 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_34_345 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_36_346 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_38_347 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_40_348 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_42_349 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_44_350 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_46_351 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_48_352 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_50_353 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_52_354 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_54_355 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_56_356 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_58_357 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_60_358 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_62_359 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_64_360 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_66_361 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_68_362 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_70_363 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_72_364 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_74_365 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_76_366 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_78_367 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_80_368 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_82_369 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_84_370 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_86_371 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_88_372 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_90_373 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_92_374 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_94_375 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_96_376 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_98_377 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_100_378 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_102_379 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_104_380 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_106_381 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_108_382 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_110_383 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_112_384 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_114_385 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_116_386 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_118_387 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_120_388 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_122_389 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_124_390 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_126_391 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_128_392 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_130_393 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_132_394 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_134_395 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_136_396 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_138_397 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_140_398 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_142_399 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_144_400 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_146_401 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_148_402 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_150_403 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_152_404 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_154_405 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_156_406 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_158_407 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_160_408 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_162_409 ();
 TAPCELL_X1 TAP_TAPCELL_ROW_163_410 ();
 BUF_X2 wire1 (.A(_00081_),
    .Z(net9));
 BUF_X4 max_cap2 (.A(_14893_),
    .Z(net10));
 BUF_X4 wire3 (.A(_04306_),
    .Z(net11));
 BUF_X4 wire4 (.A(_04302_),
    .Z(net17));
 BUF_X2 input1 (.A(key[0]),
    .Z(net19));
 BUF_X1 input2 (.A(key[100]),
    .Z(net20));
 CLKBUF_X2 input3 (.A(key[101]),
    .Z(net21));
 BUF_X1 input4 (.A(key[102]),
    .Z(net22));
 BUF_X1 input5 (.A(key[103]),
    .Z(net23));
 BUF_X1 input6 (.A(key[104]),
    .Z(net24));
 BUF_X1 input7 (.A(key[105]),
    .Z(net25));
 BUF_X1 input8 (.A(key[106]),
    .Z(net26));
 CLKBUF_X2 input9 (.A(key[107]),
    .Z(net30));
 BUF_X2 input10 (.A(key[108]),
    .Z(net31));
 BUF_X1 input11 (.A(key[109]),
    .Z(net33));
 CLKBUF_X2 input12 (.A(key[10]),
    .Z(net34));
 BUF_X2 input13 (.A(key[110]),
    .Z(net35));
 BUF_X1 input14 (.A(key[111]),
    .Z(net38));
 CLKBUF_X2 input15 (.A(key[112]),
    .Z(net40));
 BUF_X1 input16 (.A(key[113]),
    .Z(net41));
 CLKBUF_X2 input17 (.A(key[114]),
    .Z(net44));
 CLKBUF_X2 input18 (.A(key[115]),
    .Z(net45));
 BUF_X1 input19 (.A(key[116]),
    .Z(net46));
 BUF_X1 input20 (.A(key[117]),
    .Z(net47));
 CLKBUF_X2 input21 (.A(key[118]),
    .Z(net48));
 BUF_X1 input22 (.A(key[119]),
    .Z(net50));
 BUF_X2 input23 (.A(key[11]),
    .Z(net52));
 BUF_X2 input24 (.A(key[120]),
    .Z(net53));
 BUF_X2 input25 (.A(key[121]),
    .Z(net54));
 BUF_X2 input26 (.A(key[122]),
    .Z(net55));
 BUF_X2 input27 (.A(key[123]),
    .Z(net56));
 BUF_X2 input28 (.A(key[124]),
    .Z(net58));
 BUF_X2 input29 (.A(key[125]),
    .Z(net59));
 BUF_X2 input30 (.A(key[126]),
    .Z(net60));
 BUF_X2 input31 (.A(key[127]),
    .Z(net61));
 BUF_X1 input32 (.A(key[12]),
    .Z(net62));
 CLKBUF_X2 input33 (.A(key[13]),
    .Z(net63));
 CLKBUF_X2 input34 (.A(key[14]),
    .Z(net67));
 BUF_X2 input35 (.A(key[15]),
    .Z(net68));
 BUF_X1 input36 (.A(key[16]),
    .Z(net69));
 CLKBUF_X2 input37 (.A(key[17]),
    .Z(net70));
 CLKBUF_X2 input38 (.A(key[18]),
    .Z(net71));
 BUF_X1 input39 (.A(key[19]),
    .Z(net72));
 BUF_X2 input40 (.A(key[1]),
    .Z(net73));
 CLKBUF_X2 input41 (.A(key[20]),
    .Z(net74));
 CLKBUF_X2 input42 (.A(key[21]),
    .Z(net75));
 BUF_X2 input43 (.A(key[22]),
    .Z(net77));
 BUF_X1 input44 (.A(key[23]),
    .Z(net78));
 BUF_X1 input45 (.A(key[24]),
    .Z(net79));
 BUF_X2 input46 (.A(key[25]),
    .Z(net80));
 BUF_X2 input47 (.A(key[26]),
    .Z(net81));
 BUF_X2 input48 (.A(key[28]),
    .Z(net82));
 BUF_X1 input49 (.A(key[29]),
    .Z(net83));
 BUF_X1 input50 (.A(key[2]),
    .Z(net84));
 BUF_X1 input51 (.A(key[30]),
    .Z(net85));
 BUF_X2 input52 (.A(key[31]),
    .Z(net86));
 BUF_X2 input53 (.A(key[32]),
    .Z(net87));
 BUF_X1 input54 (.A(key[33]),
    .Z(net88));
 BUF_X1 input55 (.A(key[34]),
    .Z(net89));
 BUF_X1 input56 (.A(key[35]),
    .Z(net90));
 BUF_X1 input57 (.A(key[36]),
    .Z(net91));
 CLKBUF_X2 input58 (.A(key[37]),
    .Z(net92));
 BUF_X1 input59 (.A(key[38]),
    .Z(net104));
 BUF_X2 input60 (.A(key[39]),
    .Z(net115));
 BUF_X2 input61 (.A(key[3]),
    .Z(net116));
 BUF_X2 input62 (.A(key[40]),
    .Z(net117));
 CLKBUF_X2 input63 (.A(key[41]),
    .Z(net118));
 BUF_X2 input64 (.A(key[42]),
    .Z(net119));
 BUF_X1 input65 (.A(key[43]),
    .Z(net120));
 BUF_X1 input66 (.A(key[44]),
    .Z(net121));
 BUF_X1 input67 (.A(key[45]),
    .Z(net127));
 BUF_X1 input68 (.A(key[46]),
    .Z(net128));
 BUF_X1 input69 (.A(key[47]),
    .Z(net129));
 BUF_X1 input70 (.A(key[48]),
    .Z(net130));
 BUF_X1 input71 (.A(key[49]),
    .Z(net131));
 BUF_X1 input72 (.A(key[4]),
    .Z(net132));
 BUF_X2 input73 (.A(key[50]),
    .Z(net134));
 BUF_X2 input74 (.A(key[51]),
    .Z(net135));
 BUF_X1 input75 (.A(key[52]),
    .Z(net136));
 BUF_X1 input76 (.A(key[53]),
    .Z(net137));
 BUF_X1 input77 (.A(key[54]),
    .Z(net142));
 BUF_X2 input78 (.A(key[55]),
    .Z(net147));
 BUF_X1 input79 (.A(key[56]),
    .Z(net148));
 BUF_X1 input80 (.A(key[57]),
    .Z(net150));
 BUF_X1 input81 (.A(key[58]),
    .Z(net151));
 BUF_X1 input82 (.A(key[59]),
    .Z(net158));
 BUF_X1 input83 (.A(key[5]),
    .Z(net163));
 BUF_X1 input84 (.A(key[60]),
    .Z(net164));
 BUF_X1 input85 (.A(key[61]),
    .Z(net167));
 BUF_X1 input86 (.A(key[62]),
    .Z(net168));
 BUF_X1 input87 (.A(key[63]),
    .Z(net169));
 BUF_X1 input88 (.A(key[64]),
    .Z(net170));
 BUF_X1 input89 (.A(key[65]),
    .Z(net172));
 BUF_X1 input90 (.A(key[66]),
    .Z(net179));
 BUF_X1 input91 (.A(key[67]),
    .Z(net180));
 BUF_X1 input92 (.A(key[68]),
    .Z(net181));
 CLKBUF_X2 input93 (.A(key[69]),
    .Z(net182));
 BUF_X1 input94 (.A(key[6]),
    .Z(net183));
 BUF_X1 input95 (.A(key[70]),
    .Z(net184));
 BUF_X2 input96 (.A(key[71]),
    .Z(net185));
 BUF_X2 input97 (.A(key[72]),
    .Z(net186));
 BUF_X2 input98 (.A(key[73]),
    .Z(net190));
 BUF_X2 input99 (.A(key[74]),
    .Z(net191));
 CLKBUF_X2 input100 (.A(key[75]),
    .Z(net192));
 BUF_X2 input101 (.A(key[76]),
    .Z(net193));
 BUF_X2 input102 (.A(key[77]),
    .Z(net194));
 CLKBUF_X2 input103 (.A(key[78]),
    .Z(net198));
 BUF_X1 input104 (.A(key[79]),
    .Z(net199));
 BUF_X2 input105 (.A(key[7]),
    .Z(net201));
 CLKBUF_X2 input106 (.A(key[80]),
    .Z(net204));
 BUF_X1 input107 (.A(key[81]),
    .Z(net205));
 BUF_X2 input108 (.A(key[82]),
    .Z(net206));
 BUF_X2 input109 (.A(key[83]),
    .Z(net207));
 BUF_X1 input110 (.A(key[84]),
    .Z(net208));
 BUF_X1 input111 (.A(key[85]),
    .Z(net209));
 BUF_X2 input112 (.A(key[86]),
    .Z(net210));
 BUF_X2 input113 (.A(key[87]),
    .Z(net211));
 BUF_X1 input114 (.A(key[88]),
    .Z(net212));
 BUF_X1 input115 (.A(key[89]),
    .Z(net213));
 CLKBUF_X3 input116 (.A(key[8]),
    .Z(net214));
 BUF_X1 input117 (.A(key[90]),
    .Z(net215));
 BUF_X1 input118 (.A(key[91]),
    .Z(net216));
 BUF_X1 input119 (.A(key[92]),
    .Z(net217));
 BUF_X1 input120 (.A(key[93]),
    .Z(net218));
 BUF_X1 input121 (.A(key[94]),
    .Z(net219));
 BUF_X1 input122 (.A(key[95]),
    .Z(net220));
 BUF_X1 input123 (.A(key[96]),
    .Z(net221));
 BUF_X1 input124 (.A(key[97]),
    .Z(net222));
 BUF_X1 input125 (.A(key[98]),
    .Z(net223));
 BUF_X1 input126 (.A(key[99]),
    .Z(net224));
 BUF_X1 input127 (.A(key[9]),
    .Z(net225));
 CLKBUF_X3 input128 (.A(ld),
    .Z(net226));
 CLKBUF_X2 input129 (.A(rst),
    .Z(net227));
 BUF_X1 input130 (.A(text_in[0]),
    .Z(net228));
 BUF_X1 input131 (.A(text_in[100]),
    .Z(net229));
 CLKBUF_X2 input132 (.A(text_in[101]),
    .Z(net230));
 CLKBUF_X2 input133 (.A(text_in[102]),
    .Z(net231));
 CLKBUF_X2 input134 (.A(text_in[103]),
    .Z(net232));
 BUF_X1 input135 (.A(text_in[104]),
    .Z(net233));
 BUF_X1 input136 (.A(text_in[105]),
    .Z(net234));
 BUF_X2 input137 (.A(text_in[106]),
    .Z(net235));
 BUF_X1 input138 (.A(text_in[107]),
    .Z(net236));
 BUF_X1 input139 (.A(text_in[108]),
    .Z(net237));
 BUF_X1 input140 (.A(text_in[109]),
    .Z(net238));
 BUF_X1 input141 (.A(text_in[10]),
    .Z(net239));
 BUF_X1 input142 (.A(text_in[110]),
    .Z(net240));
 BUF_X1 input143 (.A(text_in[111]),
    .Z(net241));
 BUF_X1 input144 (.A(text_in[112]),
    .Z(net242));
 BUF_X1 input145 (.A(text_in[113]),
    .Z(net243));
 BUF_X1 input146 (.A(text_in[114]),
    .Z(net244));
 BUF_X1 input147 (.A(text_in[115]),
    .Z(net245));
 BUF_X1 input148 (.A(text_in[116]),
    .Z(net246));
 BUF_X1 input149 (.A(text_in[117]),
    .Z(net247));
 BUF_X1 input150 (.A(text_in[118]),
    .Z(net248));
 BUF_X1 input151 (.A(text_in[119]),
    .Z(net249));
 BUF_X1 input152 (.A(text_in[11]),
    .Z(net250));
 BUF_X1 input153 (.A(text_in[120]),
    .Z(net251));
 BUF_X2 input154 (.A(text_in[121]),
    .Z(net252));
 BUF_X1 input155 (.A(text_in[122]),
    .Z(net253));
 BUF_X1 input156 (.A(text_in[123]),
    .Z(net254));
 BUF_X1 input157 (.A(text_in[124]),
    .Z(net255));
 BUF_X1 input158 (.A(text_in[125]),
    .Z(net256));
 BUF_X1 input159 (.A(text_in[126]),
    .Z(net257));
 BUF_X1 input160 (.A(text_in[127]),
    .Z(net258));
 BUF_X1 input161 (.A(text_in[12]),
    .Z(net259));
 BUF_X1 input162 (.A(text_in[13]),
    .Z(net260));
 BUF_X1 input163 (.A(text_in[14]),
    .Z(net261));
 BUF_X1 input164 (.A(text_in[15]),
    .Z(net262));
 BUF_X1 input165 (.A(text_in[16]),
    .Z(net263));
 BUF_X1 input166 (.A(text_in[17]),
    .Z(net264));
 BUF_X1 input167 (.A(text_in[18]),
    .Z(net265));
 BUF_X1 input168 (.A(text_in[19]),
    .Z(net266));
 BUF_X1 input169 (.A(text_in[1]),
    .Z(net267));
 BUF_X1 input170 (.A(text_in[20]),
    .Z(net268));
 BUF_X1 input171 (.A(text_in[21]),
    .Z(net269));
 BUF_X1 input172 (.A(text_in[22]),
    .Z(net270));
 BUF_X1 input173 (.A(text_in[23]),
    .Z(net271));
 CLKBUF_X2 input174 (.A(text_in[24]),
    .Z(net272));
 BUF_X1 input175 (.A(text_in[25]),
    .Z(net273));
 BUF_X1 input176 (.A(text_in[26]),
    .Z(net274));
 BUF_X1 input177 (.A(text_in[27]),
    .Z(net275));
 BUF_X1 input178 (.A(text_in[28]),
    .Z(net276));
 BUF_X1 input179 (.A(text_in[29]),
    .Z(net277));
 BUF_X1 input180 (.A(text_in[2]),
    .Z(net278));
 BUF_X1 input181 (.A(text_in[30]),
    .Z(net279));
 BUF_X1 input182 (.A(text_in[31]),
    .Z(net280));
 BUF_X1 input183 (.A(text_in[32]),
    .Z(net281));
 BUF_X1 input184 (.A(text_in[33]),
    .Z(net282));
 CLKBUF_X2 input185 (.A(text_in[34]),
    .Z(net283));
 BUF_X1 input186 (.A(text_in[35]),
    .Z(net284));
 BUF_X1 input187 (.A(text_in[36]),
    .Z(net285));
 BUF_X1 input188 (.A(text_in[37]),
    .Z(net286));
 CLKBUF_X2 input189 (.A(text_in[38]),
    .Z(net287));
 BUF_X1 input190 (.A(text_in[39]),
    .Z(net288));
 BUF_X1 input191 (.A(text_in[3]),
    .Z(net289));
 BUF_X1 input192 (.A(text_in[40]),
    .Z(net290));
 BUF_X1 input193 (.A(text_in[41]),
    .Z(net291));
 BUF_X1 input194 (.A(text_in[42]),
    .Z(net292));
 BUF_X1 input195 (.A(text_in[43]),
    .Z(net293));
 BUF_X1 input196 (.A(text_in[44]),
    .Z(net294));
 CLKBUF_X2 input197 (.A(text_in[45]),
    .Z(net295));
 BUF_X1 input198 (.A(text_in[46]),
    .Z(net296));
 BUF_X1 input199 (.A(text_in[47]),
    .Z(net297));
 BUF_X1 input200 (.A(text_in[48]),
    .Z(net298));
 BUF_X1 input201 (.A(text_in[49]),
    .Z(net299));
 BUF_X1 input202 (.A(text_in[4]),
    .Z(net300));
 BUF_X1 input203 (.A(text_in[50]),
    .Z(net301));
 BUF_X1 input204 (.A(text_in[51]),
    .Z(net302));
 BUF_X1 input205 (.A(text_in[52]),
    .Z(net303));
 BUF_X1 input206 (.A(text_in[53]),
    .Z(net304));
 BUF_X1 input207 (.A(text_in[54]),
    .Z(net305));
 BUF_X1 input208 (.A(text_in[55]),
    .Z(net306));
 BUF_X1 input209 (.A(text_in[56]),
    .Z(net307));
 BUF_X1 input210 (.A(text_in[57]),
    .Z(net308));
 BUF_X1 input211 (.A(text_in[58]),
    .Z(net309));
 BUF_X1 input212 (.A(text_in[59]),
    .Z(net310));
 BUF_X1 input213 (.A(text_in[5]),
    .Z(net311));
 BUF_X1 input214 (.A(text_in[60]),
    .Z(net312));
 BUF_X1 input215 (.A(text_in[61]),
    .Z(net313));
 BUF_X1 input216 (.A(text_in[62]),
    .Z(net314));
 BUF_X1 input217 (.A(text_in[63]),
    .Z(net315));
 BUF_X1 input218 (.A(text_in[64]),
    .Z(net316));
 BUF_X1 input219 (.A(text_in[65]),
    .Z(net317));
 BUF_X1 input220 (.A(text_in[66]),
    .Z(net318));
 BUF_X1 input221 (.A(text_in[67]),
    .Z(net319));
 BUF_X1 input222 (.A(text_in[68]),
    .Z(net320));
 BUF_X1 input223 (.A(text_in[69]),
    .Z(net321));
 BUF_X1 input224 (.A(text_in[6]),
    .Z(net322));
 BUF_X1 input225 (.A(text_in[70]),
    .Z(net323));
 BUF_X1 input226 (.A(text_in[71]),
    .Z(net324));
 CLKBUF_X2 input227 (.A(text_in[72]),
    .Z(net325));
 BUF_X1 input228 (.A(text_in[73]),
    .Z(net326));
 BUF_X1 input229 (.A(text_in[74]),
    .Z(net327));
 BUF_X1 input230 (.A(text_in[75]),
    .Z(net328));
 BUF_X1 input231 (.A(text_in[76]),
    .Z(net329));
 BUF_X2 input232 (.A(text_in[77]),
    .Z(net330));
 CLKBUF_X2 input233 (.A(text_in[78]),
    .Z(net331));
 BUF_X1 input234 (.A(text_in[79]),
    .Z(net332));
 BUF_X1 input235 (.A(text_in[7]),
    .Z(net333));
 CLKBUF_X2 input236 (.A(text_in[80]),
    .Z(net334));
 CLKBUF_X2 input237 (.A(text_in[81]),
    .Z(net335));
 CLKBUF_X2 input238 (.A(text_in[82]),
    .Z(net336));
 CLKBUF_X2 input239 (.A(text_in[83]),
    .Z(net337));
 BUF_X1 input240 (.A(text_in[84]),
    .Z(net338));
 BUF_X1 input241 (.A(text_in[85]),
    .Z(net339));
 BUF_X1 input242 (.A(text_in[86]),
    .Z(net340));
 BUF_X1 input243 (.A(text_in[87]),
    .Z(net341));
 BUF_X1 input244 (.A(text_in[88]),
    .Z(net342));
 BUF_X1 input245 (.A(text_in[89]),
    .Z(net343));
 CLKBUF_X2 input246 (.A(text_in[8]),
    .Z(net344));
 BUF_X1 input247 (.A(text_in[90]),
    .Z(net345));
 BUF_X1 input248 (.A(text_in[91]),
    .Z(net346));
 BUF_X1 input249 (.A(text_in[92]),
    .Z(net347));
 BUF_X1 input250 (.A(text_in[93]),
    .Z(net348));
 BUF_X1 input251 (.A(text_in[94]),
    .Z(net349));
 BUF_X1 input252 (.A(text_in[95]),
    .Z(net350));
 BUF_X2 input253 (.A(text_in[96]),
    .Z(net351));
 BUF_X1 input254 (.A(text_in[97]),
    .Z(net352));
 BUF_X1 input255 (.A(text_in[98]),
    .Z(net353));
 BUF_X1 input256 (.A(text_in[99]),
    .Z(net354));
 BUF_X1 input257 (.A(text_in[9]),
    .Z(net355));
 BUF_X1 output258 (.A(net356),
    .Z(done));
 BUF_X1 output259 (.A(net357),
    .Z(text_out[0]));
 BUF_X1 output260 (.A(net358),
    .Z(text_out[100]));
 BUF_X1 output261 (.A(net359),
    .Z(text_out[101]));
 BUF_X1 output262 (.A(net360),
    .Z(text_out[102]));
 BUF_X1 output263 (.A(net361),
    .Z(text_out[103]));
 BUF_X1 output264 (.A(net362),
    .Z(text_out[104]));
 BUF_X1 output265 (.A(net363),
    .Z(text_out[105]));
 BUF_X1 output266 (.A(net364),
    .Z(text_out[106]));
 BUF_X1 output267 (.A(net365),
    .Z(text_out[107]));
 BUF_X1 output268 (.A(net366),
    .Z(text_out[108]));
 BUF_X1 output269 (.A(net367),
    .Z(text_out[109]));
 BUF_X1 output270 (.A(net368),
    .Z(text_out[10]));
 BUF_X1 output271 (.A(net369),
    .Z(text_out[110]));
 BUF_X1 output272 (.A(net370),
    .Z(text_out[111]));
 BUF_X1 output273 (.A(net371),
    .Z(text_out[112]));
 BUF_X1 output274 (.A(net372),
    .Z(text_out[113]));
 BUF_X1 output275 (.A(net373),
    .Z(text_out[114]));
 BUF_X1 output276 (.A(net374),
    .Z(text_out[115]));
 BUF_X1 output277 (.A(net375),
    .Z(text_out[116]));
 BUF_X1 output278 (.A(net376),
    .Z(text_out[117]));
 BUF_X1 output279 (.A(net377),
    .Z(text_out[118]));
 BUF_X1 output280 (.A(net378),
    .Z(text_out[119]));
 BUF_X1 output281 (.A(net379),
    .Z(text_out[11]));
 BUF_X1 output282 (.A(net380),
    .Z(text_out[120]));
 BUF_X1 output283 (.A(net381),
    .Z(text_out[121]));
 BUF_X1 output284 (.A(net382),
    .Z(text_out[122]));
 BUF_X1 output285 (.A(net383),
    .Z(text_out[123]));
 BUF_X1 output286 (.A(net384),
    .Z(text_out[124]));
 BUF_X1 output287 (.A(net385),
    .Z(text_out[125]));
 BUF_X1 output288 (.A(net386),
    .Z(text_out[126]));
 BUF_X1 output289 (.A(net387),
    .Z(text_out[127]));
 BUF_X1 output290 (.A(net388),
    .Z(text_out[12]));
 BUF_X1 output291 (.A(net389),
    .Z(text_out[13]));
 BUF_X1 output292 (.A(net390),
    .Z(text_out[14]));
 BUF_X1 output293 (.A(net391),
    .Z(text_out[15]));
 BUF_X1 output294 (.A(net392),
    .Z(text_out[16]));
 BUF_X1 output295 (.A(net393),
    .Z(text_out[17]));
 BUF_X1 output296 (.A(net394),
    .Z(text_out[18]));
 BUF_X1 output297 (.A(net395),
    .Z(text_out[19]));
 BUF_X1 output298 (.A(net396),
    .Z(text_out[1]));
 BUF_X1 output299 (.A(net397),
    .Z(text_out[20]));
 BUF_X1 output300 (.A(net398),
    .Z(text_out[21]));
 BUF_X1 output301 (.A(net399),
    .Z(text_out[22]));
 BUF_X1 output302 (.A(net400),
    .Z(text_out[23]));
 BUF_X1 output303 (.A(net401),
    .Z(text_out[24]));
 BUF_X1 output304 (.A(net402),
    .Z(text_out[25]));
 BUF_X1 output305 (.A(net403),
    .Z(text_out[26]));
 BUF_X1 output306 (.A(net404),
    .Z(text_out[27]));
 BUF_X1 output307 (.A(net405),
    .Z(text_out[28]));
 BUF_X1 output308 (.A(net406),
    .Z(text_out[29]));
 BUF_X1 output309 (.A(net407),
    .Z(text_out[2]));
 BUF_X1 output310 (.A(net408),
    .Z(text_out[30]));
 BUF_X1 output311 (.A(net409),
    .Z(text_out[31]));
 BUF_X1 output312 (.A(net410),
    .Z(text_out[32]));
 BUF_X1 output313 (.A(net411),
    .Z(text_out[33]));
 BUF_X1 output314 (.A(net412),
    .Z(text_out[34]));
 BUF_X1 output315 (.A(net413),
    .Z(text_out[35]));
 BUF_X1 output316 (.A(net414),
    .Z(text_out[36]));
 BUF_X1 output317 (.A(net415),
    .Z(text_out[37]));
 BUF_X1 output318 (.A(net416),
    .Z(text_out[38]));
 BUF_X1 output319 (.A(net417),
    .Z(text_out[39]));
 BUF_X1 output320 (.A(net418),
    .Z(text_out[3]));
 BUF_X1 output321 (.A(net419),
    .Z(text_out[40]));
 BUF_X1 output322 (.A(net420),
    .Z(text_out[41]));
 BUF_X1 output323 (.A(net421),
    .Z(text_out[42]));
 BUF_X1 output324 (.A(net422),
    .Z(text_out[43]));
 BUF_X1 output325 (.A(net423),
    .Z(text_out[44]));
 BUF_X1 output326 (.A(net424),
    .Z(text_out[45]));
 BUF_X1 output327 (.A(net425),
    .Z(text_out[46]));
 BUF_X1 output328 (.A(net426),
    .Z(text_out[47]));
 BUF_X1 output329 (.A(net427),
    .Z(text_out[48]));
 BUF_X1 output330 (.A(net428),
    .Z(text_out[49]));
 BUF_X1 output331 (.A(net429),
    .Z(text_out[4]));
 BUF_X1 output332 (.A(net430),
    .Z(text_out[50]));
 BUF_X1 output333 (.A(net431),
    .Z(text_out[51]));
 BUF_X1 output334 (.A(net432),
    .Z(text_out[52]));
 BUF_X1 output335 (.A(net433),
    .Z(text_out[53]));
 BUF_X1 output336 (.A(net434),
    .Z(text_out[54]));
 BUF_X1 output337 (.A(net435),
    .Z(text_out[55]));
 BUF_X1 output338 (.A(net436),
    .Z(text_out[56]));
 BUF_X1 output339 (.A(net437),
    .Z(text_out[57]));
 BUF_X1 output340 (.A(net438),
    .Z(text_out[58]));
 BUF_X1 output341 (.A(net439),
    .Z(text_out[59]));
 BUF_X1 output342 (.A(net440),
    .Z(text_out[5]));
 BUF_X1 output343 (.A(net441),
    .Z(text_out[60]));
 BUF_X1 output344 (.A(net442),
    .Z(text_out[61]));
 BUF_X1 output345 (.A(net443),
    .Z(text_out[62]));
 BUF_X1 output346 (.A(net444),
    .Z(text_out[63]));
 BUF_X1 output347 (.A(net445),
    .Z(text_out[64]));
 BUF_X1 output348 (.A(net446),
    .Z(text_out[65]));
 BUF_X1 output349 (.A(net447),
    .Z(text_out[66]));
 BUF_X1 output350 (.A(net448),
    .Z(text_out[67]));
 BUF_X1 output351 (.A(net449),
    .Z(text_out[68]));
 BUF_X1 output352 (.A(net450),
    .Z(text_out[69]));
 BUF_X1 output353 (.A(net451),
    .Z(text_out[6]));
 BUF_X1 output354 (.A(net452),
    .Z(text_out[70]));
 BUF_X1 output355 (.A(net453),
    .Z(text_out[71]));
 BUF_X1 output356 (.A(net454),
    .Z(text_out[72]));
 BUF_X1 output357 (.A(net455),
    .Z(text_out[73]));
 BUF_X1 output358 (.A(net456),
    .Z(text_out[74]));
 BUF_X1 output359 (.A(net457),
    .Z(text_out[75]));
 BUF_X1 output360 (.A(net458),
    .Z(text_out[76]));
 BUF_X1 output361 (.A(net459),
    .Z(text_out[77]));
 BUF_X1 output362 (.A(net460),
    .Z(text_out[78]));
 BUF_X1 output363 (.A(net461),
    .Z(text_out[79]));
 BUF_X1 output364 (.A(net462),
    .Z(text_out[7]));
 BUF_X1 output365 (.A(net463),
    .Z(text_out[80]));
 BUF_X1 output366 (.A(net464),
    .Z(text_out[81]));
 BUF_X1 output367 (.A(net465),
    .Z(text_out[82]));
 BUF_X1 output368 (.A(net466),
    .Z(text_out[83]));
 BUF_X1 output369 (.A(net467),
    .Z(text_out[84]));
 BUF_X1 output370 (.A(net468),
    .Z(text_out[85]));
 BUF_X1 output371 (.A(net469),
    .Z(text_out[86]));
 BUF_X1 output372 (.A(net470),
    .Z(text_out[87]));
 BUF_X1 output373 (.A(net471),
    .Z(text_out[88]));
 BUF_X1 output374 (.A(net472),
    .Z(text_out[89]));
 BUF_X1 output375 (.A(net473),
    .Z(text_out[8]));
 BUF_X1 output376 (.A(net474),
    .Z(text_out[90]));
 BUF_X1 output377 (.A(net475),
    .Z(text_out[91]));
 BUF_X1 output378 (.A(net476),
    .Z(text_out[92]));
 BUF_X1 output379 (.A(net477),
    .Z(text_out[93]));
 BUF_X1 output380 (.A(net478),
    .Z(text_out[94]));
 BUF_X1 output381 (.A(net479),
    .Z(text_out[95]));
 BUF_X1 output382 (.A(net480),
    .Z(text_out[96]));
 BUF_X1 output383 (.A(net481),
    .Z(text_out[97]));
 BUF_X1 output384 (.A(net482),
    .Z(text_out[98]));
 BUF_X1 output385 (.A(net483),
    .Z(text_out[99]));
 BUF_X1 output386 (.A(net484),
    .Z(text_out[9]));
 CLKBUF_X3 clkbuf_leaf_0_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_0_clk));
 CLKBUF_X3 clkbuf_leaf_1_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_1_clk));
 CLKBUF_X3 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_2_clk));
 CLKBUF_X3 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_3_clk));
 CLKBUF_X3 clkbuf_leaf_4_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_4_clk));
 CLKBUF_X3 clkbuf_leaf_5_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_5_clk));
 CLKBUF_X3 clkbuf_leaf_6_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_6_clk));
 CLKBUF_X3 clkbuf_leaf_7_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_7_clk));
 CLKBUF_X3 clkbuf_leaf_8_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_8_clk));
 CLKBUF_X3 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_9_clk));
 CLKBUF_X3 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_10_clk));
 CLKBUF_X3 clkbuf_leaf_11_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_11_clk));
 CLKBUF_X3 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_12_clk));
 CLKBUF_X3 clkbuf_leaf_13_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_13_clk));
 CLKBUF_X3 clkbuf_leaf_14_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_14_clk));
 CLKBUF_X3 clkbuf_leaf_15_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_15_clk));
 CLKBUF_X3 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_16_clk));
 CLKBUF_X3 clkbuf_leaf_17_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_17_clk));
 CLKBUF_X3 clkbuf_leaf_18_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_18_clk));
 CLKBUF_X3 clkbuf_leaf_19_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_19_clk));
 CLKBUF_X3 clkbuf_leaf_20_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_20_clk));
 CLKBUF_X3 clkbuf_leaf_21_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_21_clk));
 CLKBUF_X3 clkbuf_leaf_22_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_22_clk));
 CLKBUF_X3 clkbuf_leaf_23_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_23_clk));
 CLKBUF_X3 clkbuf_leaf_24_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_24_clk));
 CLKBUF_X3 clkbuf_leaf_25_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_25_clk));
 CLKBUF_X3 clkbuf_leaf_26_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_26_clk));
 CLKBUF_X3 clkbuf_leaf_27_clk (.A(clknet_3_3__leaf_clk),
    .Z(clknet_leaf_27_clk));
 CLKBUF_X3 clkbuf_leaf_28_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_28_clk));
 CLKBUF_X3 clkbuf_leaf_29_clk (.A(clknet_3_2__leaf_clk),
    .Z(clknet_leaf_29_clk));
 CLKBUF_X3 clkbuf_leaf_30_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_30_clk));
 CLKBUF_X3 clkbuf_leaf_31_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_31_clk));
 CLKBUF_X3 clkbuf_leaf_32_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_32_clk));
 CLKBUF_X3 clkbuf_leaf_33_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_33_clk));
 CLKBUF_X3 clkbuf_leaf_34_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_34_clk));
 CLKBUF_X3 clkbuf_leaf_35_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_35_clk));
 CLKBUF_X3 clkbuf_leaf_36_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_36_clk));
 CLKBUF_X3 clkbuf_leaf_37_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_37_clk));
 CLKBUF_X3 clkbuf_leaf_38_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_38_clk));
 CLKBUF_X3 clkbuf_leaf_39_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_39_clk));
 CLKBUF_X3 clkbuf_leaf_40_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_40_clk));
 CLKBUF_X3 clkbuf_leaf_41_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_41_clk));
 CLKBUF_X3 clkbuf_leaf_42_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_42_clk));
 CLKBUF_X3 clkbuf_leaf_43_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_43_clk));
 CLKBUF_X3 clkbuf_leaf_44_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_44_clk));
 CLKBUF_X3 clkbuf_leaf_45_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_45_clk));
 CLKBUF_X3 clkbuf_leaf_46_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_46_clk));
 CLKBUF_X3 clkbuf_leaf_47_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_47_clk));
 CLKBUF_X3 clkbuf_leaf_48_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_48_clk));
 CLKBUF_X3 clkbuf_leaf_49_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_49_clk));
 CLKBUF_X3 clkbuf_leaf_50_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_50_clk));
 CLKBUF_X3 clkbuf_leaf_51_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_51_clk));
 CLKBUF_X3 clkbuf_leaf_52_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_52_clk));
 CLKBUF_X3 clkbuf_leaf_53_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_53_clk));
 CLKBUF_X3 clkbuf_leaf_54_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_54_clk));
 CLKBUF_X3 clkbuf_leaf_55_clk (.A(clknet_3_7__leaf_clk),
    .Z(clknet_leaf_55_clk));
 CLKBUF_X3 clkbuf_leaf_56_clk (.A(clknet_3_6__leaf_clk),
    .Z(clknet_leaf_56_clk));
 CLKBUF_X3 clkbuf_leaf_57_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_57_clk));
 CLKBUF_X3 clkbuf_leaf_58_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_58_clk));
 CLKBUF_X3 clkbuf_leaf_59_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_59_clk));
 CLKBUF_X3 clkbuf_leaf_60_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_60_clk));
 CLKBUF_X3 clkbuf_leaf_61_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_61_clk));
 CLKBUF_X3 clkbuf_leaf_62_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_62_clk));
 CLKBUF_X3 clkbuf_leaf_63_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_63_clk));
 CLKBUF_X3 clkbuf_leaf_64_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_64_clk));
 CLKBUF_X3 clkbuf_leaf_65_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_65_clk));
 CLKBUF_X3 clkbuf_leaf_66_clk (.A(clknet_3_5__leaf_clk),
    .Z(clknet_leaf_66_clk));
 CLKBUF_X3 clkbuf_leaf_67_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_67_clk));
 CLKBUF_X3 clkbuf_leaf_68_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_68_clk));
 CLKBUF_X3 clkbuf_leaf_69_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_69_clk));
 CLKBUF_X3 clkbuf_leaf_70_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_70_clk));
 CLKBUF_X3 clkbuf_leaf_71_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_71_clk));
 CLKBUF_X3 clkbuf_leaf_72_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_72_clk));
 CLKBUF_X3 clkbuf_leaf_73_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_73_clk));
 CLKBUF_X3 clkbuf_leaf_74_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_74_clk));
 CLKBUF_X3 clkbuf_leaf_75_clk (.A(clknet_3_4__leaf_clk),
    .Z(clknet_leaf_75_clk));
 CLKBUF_X3 clkbuf_leaf_76_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_76_clk));
 CLKBUF_X3 clkbuf_leaf_77_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_77_clk));
 CLKBUF_X3 clkbuf_leaf_78_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_78_clk));
 CLKBUF_X3 clkbuf_leaf_79_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_79_clk));
 CLKBUF_X3 clkbuf_leaf_80_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_80_clk));
 CLKBUF_X3 clkbuf_leaf_81_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_81_clk));
 CLKBUF_X3 clkbuf_leaf_82_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_82_clk));
 CLKBUF_X3 clkbuf_leaf_83_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_83_clk));
 CLKBUF_X3 clkbuf_leaf_84_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_84_clk));
 CLKBUF_X3 clkbuf_leaf_85_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_85_clk));
 CLKBUF_X3 clkbuf_leaf_86_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_86_clk));
 CLKBUF_X3 clkbuf_leaf_87_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_87_clk));
 CLKBUF_X3 clkbuf_leaf_88_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_88_clk));
 CLKBUF_X3 clkbuf_leaf_89_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_89_clk));
 CLKBUF_X3 clkbuf_leaf_90_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_90_clk));
 CLKBUF_X3 clkbuf_leaf_91_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_91_clk));
 CLKBUF_X3 clkbuf_leaf_92_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_92_clk));
 CLKBUF_X3 clkbuf_leaf_93_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_93_clk));
 CLKBUF_X3 clkbuf_leaf_94_clk (.A(clknet_3_1__leaf_clk),
    .Z(clknet_leaf_94_clk));
 CLKBUF_X3 clkbuf_leaf_95_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_95_clk));
 CLKBUF_X3 clkbuf_leaf_96_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_96_clk));
 CLKBUF_X3 clkbuf_leaf_97_clk (.A(clknet_3_0__leaf_clk),
    .Z(clknet_leaf_97_clk));
 CLKBUF_X3 clkbuf_0_clk (.A(clk),
    .Z(clknet_0_clk));
 CLKBUF_X3 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_0__leaf_clk));
 CLKBUF_X3 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_1__leaf_clk));
 CLKBUF_X3 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_2__leaf_clk));
 CLKBUF_X3 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_3__leaf_clk));
 CLKBUF_X3 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_4__leaf_clk));
 CLKBUF_X3 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_5__leaf_clk));
 CLKBUF_X3 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_6__leaf_clk));
 CLKBUF_X3 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .Z(clknet_3_7__leaf_clk));
 INV_X4 clkload0 (.A(clknet_3_0__leaf_clk));
 INV_X2 clkload1 (.A(clknet_3_2__leaf_clk));
 INV_X8 clkload2 (.A(clknet_3_3__leaf_clk));
 INV_X8 clkload3 (.A(clknet_3_4__leaf_clk));
 INV_X2 clkload4 (.A(clknet_3_5__leaf_clk));
 INV_X8 clkload5 (.A(clknet_3_6__leaf_clk));
 INV_X4 clkload6 (.A(clknet_3_7__leaf_clk));
 INV_X1 clkload7 (.A(clknet_leaf_2_clk));
 INV_X2 clkload8 (.A(clknet_leaf_3_clk));
 INV_X2 clkload9 (.A(clknet_leaf_6_clk));
 CLKBUF_X1 clkload10 (.A(clknet_leaf_85_clk));
 INV_X1 clkload11 (.A(clknet_leaf_86_clk));
 INV_X2 clkload12 (.A(clknet_leaf_87_clk));
 INV_X1 clkload13 (.A(clknet_leaf_88_clk));
 INV_X2 clkload14 (.A(clknet_leaf_89_clk));
 INV_X2 clkload15 (.A(clknet_leaf_95_clk));
 INV_X1 clkload16 (.A(clknet_leaf_96_clk));
 INV_X2 clkload17 (.A(clknet_leaf_97_clk));
 INV_X1 clkload18 (.A(clknet_leaf_7_clk));
 INV_X1 clkload19 (.A(clknet_leaf_8_clk));
 CLKBUF_X1 clkload20 (.A(clknet_leaf_73_clk));
 INV_X1 clkload21 (.A(clknet_leaf_74_clk));
 INV_X1 clkload22 (.A(clknet_leaf_76_clk));
 INV_X2 clkload23 (.A(clknet_leaf_77_clk));
 CLKBUF_X1 clkload24 (.A(clknet_leaf_78_clk));
 CLKBUF_X1 clkload25 (.A(clknet_leaf_79_clk));
 CLKBUF_X1 clkload26 (.A(clknet_leaf_80_clk));
 INV_X1 clkload27 (.A(clknet_leaf_81_clk));
 CLKBUF_X1 clkload28 (.A(clknet_leaf_83_clk));
 CLKBUF_X1 clkload29 (.A(clknet_leaf_84_clk));
 INV_X1 clkload30 (.A(clknet_leaf_91_clk));
 CLKBUF_X1 clkload31 (.A(clknet_leaf_92_clk));
 CLKBUF_X1 clkload32 (.A(clknet_leaf_93_clk));
 INV_X1 clkload33 (.A(clknet_leaf_94_clk));
 CLKBUF_X1 clkload34 (.A(clknet_leaf_0_clk));
 INV_X1 clkload35 (.A(clknet_leaf_1_clk));
 INV_X1 clkload36 (.A(clknet_leaf_4_clk));
 INV_X1 clkload37 (.A(clknet_leaf_5_clk));
 CLKBUF_X1 clkload38 (.A(clknet_leaf_11_clk));
 INV_X2 clkload39 (.A(clknet_leaf_12_clk));
 INV_X1 clkload40 (.A(clknet_leaf_13_clk));
 INV_X2 clkload41 (.A(clknet_leaf_16_clk));
 INV_X1 clkload42 (.A(clknet_leaf_17_clk));
 INV_X2 clkload43 (.A(clknet_leaf_18_clk));
 INV_X2 clkload44 (.A(clknet_leaf_19_clk));
 INV_X2 clkload45 (.A(clknet_leaf_20_clk));
 INV_X2 clkload46 (.A(clknet_leaf_29_clk));
 CLKBUF_X1 clkload47 (.A(clknet_leaf_10_clk));
 CLKBUF_X1 clkload48 (.A(clknet_leaf_14_clk));
 INV_X1 clkload49 (.A(clknet_leaf_15_clk));
 INV_X2 clkload50 (.A(clknet_leaf_21_clk));
 INV_X2 clkload51 (.A(clknet_leaf_22_clk));
 CLKBUF_X1 clkload52 (.A(clknet_leaf_24_clk));
 INV_X1 clkload53 (.A(clknet_leaf_25_clk));
 CLKBUF_X1 clkload54 (.A(clknet_leaf_26_clk));
 INV_X1 clkload55 (.A(clknet_leaf_27_clk));
 CLKBUF_X1 clkload56 (.A(clknet_leaf_58_clk));
 CLKBUF_X1 clkload57 (.A(clknet_leaf_60_clk));
 INV_X2 clkload58 (.A(clknet_leaf_67_clk));
 INV_X1 clkload59 (.A(clknet_leaf_68_clk));
 INV_X2 clkload60 (.A(clknet_leaf_70_clk));
 INV_X1 clkload61 (.A(clknet_leaf_71_clk));
 CLKBUF_X1 clkload62 (.A(clknet_leaf_72_clk));
 INV_X1 clkload63 (.A(clknet_leaf_75_clk));
 INV_X1 clkload64 (.A(clknet_leaf_43_clk));
 INV_X1 clkload65 (.A(clknet_leaf_44_clk));
 INV_X1 clkload66 (.A(clknet_leaf_49_clk));
 INV_X1 clkload67 (.A(clknet_leaf_57_clk));
 CLKBUF_X1 clkload68 (.A(clknet_leaf_61_clk));
 CLKBUF_X1 clkload69 (.A(clknet_leaf_62_clk));
 CLKBUF_X1 clkload70 (.A(clknet_leaf_63_clk));
 INV_X2 clkload71 (.A(clknet_leaf_64_clk));
 CLKBUF_X1 clkload72 (.A(clknet_leaf_66_clk));
 INV_X2 clkload73 (.A(clknet_leaf_28_clk));
 INV_X4 clkload74 (.A(clknet_leaf_30_clk));
 INV_X2 clkload75 (.A(clknet_leaf_31_clk));
 INV_X2 clkload76 (.A(clknet_leaf_32_clk));
 INV_X1 clkload77 (.A(clknet_leaf_34_clk));
 CLKBUF_X1 clkload78 (.A(clknet_leaf_35_clk));
 CLKBUF_X1 clkload79 (.A(clknet_leaf_36_clk));
 INV_X2 clkload80 (.A(clknet_leaf_38_clk));
 INV_X2 clkload81 (.A(clknet_leaf_56_clk));
 INV_X2 clkload82 (.A(clknet_leaf_33_clk));
 CLKBUF_X1 clkload83 (.A(clknet_leaf_39_clk));
 INV_X2 clkload84 (.A(clknet_leaf_40_clk));
 INV_X2 clkload85 (.A(clknet_leaf_42_clk));
 CLKBUF_X1 clkload86 (.A(clknet_leaf_48_clk));
 INV_X2 clkload87 (.A(clknet_leaf_50_clk));
 CLKBUF_X1 clkload88 (.A(clknet_leaf_51_clk));
 CLKBUF_X1 clkload89 (.A(clknet_leaf_52_clk));
 INV_X1 clkload90 (.A(clknet_leaf_54_clk));
 CLKBUF_X1 clkload91 (.A(clknet_leaf_55_clk));
 BUF_X4 rebuffer1 (.A(_14829_),
    .Z(net485));
 BUF_X4 rebuffer2 (.A(net485),
    .Z(net486));
 BUF_X4 rebuffer3 (.A(_13175_),
    .Z(net487));
 BUF_X1 rebuffer4 (.A(_13175_),
    .Z(net488));
 BUF_X1 rebuffer5 (.A(_14993_),
    .Z(net489));
 BUF_X1 rebuffer6 (.A(_04229_),
    .Z(net490));
 BUF_X1 rebuffer7 (.A(net490),
    .Z(net491));
 BUF_X1 rebuffer8 (.A(net490),
    .Z(net492));
 BUF_X2 rebuffer9 (.A(net490),
    .Z(net493));
 BUF_X1 rebuffer10 (.A(_13171_),
    .Z(net494));
 BUF_X2 rebuffer11 (.A(_14993_),
    .Z(net495));
 BUF_X4 rebuffer12 (.A(_09002_),
    .Z(net496));
 BUF_X1 rebuffer13 (.A(net496),
    .Z(net497));
 BUF_X2 rebuffer14 (.A(_14957_),
    .Z(net498));
 BUF_X8 rebuffer15 (.A(net498),
    .Z(net499));
 BUF_X4 rebuffer16 (.A(_14957_),
    .Z(net500));
 BUF_X8 rebuffer17 (.A(net500),
    .Z(net501));
 BUF_X1 rebuffer18 (.A(net500),
    .Z(net502));
 BUF_X4 rebuffer19 (.A(net687),
    .Z(net503));
 BUF_X2 rebuffer20 (.A(_14661_),
    .Z(net504));
 BUF_X2 rebuffer21 (.A(_06265_),
    .Z(net505));
 BUF_X2 rebuffer22 (.A(_15125_),
    .Z(net506));
 BUF_X1 rebuffer23 (.A(_04859_),
    .Z(net507));
 BUF_X1 rebuffer24 (.A(_05531_),
    .Z(net508));
 BUF_X1 rebuffer25 (.A(net883),
    .Z(net509));
 BUF_X1 rebuffer26 (.A(net509),
    .Z(net510));
 BUF_X1 rebuffer27 (.A(net509),
    .Z(net511));
 BUF_X1 rebuffer28 (.A(_03585_),
    .Z(net512));
 BUF_X2 rebuffer29 (.A(net512),
    .Z(net513));
 BUF_X1 rebuffer30 (.A(_15165_),
    .Z(net514));
 BUF_X4 rebuffer31 (.A(_15165_),
    .Z(net515));
 BUF_X1 rebuffer32 (.A(net515),
    .Z(net516));
 BUF_X4 rebuffer33 (.A(_06252_),
    .Z(net517));
 BUF_X1 rebuffer34 (.A(net517),
    .Z(net518));
 BUF_X1 rebuffer35 (.A(_00945_),
    .Z(net519));
 BUF_X1 rebuffer36 (.A(_00945_),
    .Z(net520));
 BUF_X1 rebuffer37 (.A(_10504_),
    .Z(net521));
 BUF_X2 rebuffer38 (.A(net521),
    .Z(net522));
 BUF_X1 rebuffer39 (.A(_15104_),
    .Z(net523));
 BUF_X4 rebuffer40 (.A(net789),
    .Z(net524));
 BUF_X1 rebuffer41 (.A(_08991_),
    .Z(net525));
 BUF_X1 rebuffer42 (.A(_05527_),
    .Z(net526));
 BUF_X2 rebuffer43 (.A(_05527_),
    .Z(net527));
 BUF_X1 rebuffer44 (.A(_05527_),
    .Z(net528));
 BUF_X1 rebuffer45 (.A(\sa12_sr[0] ),
    .Z(net529));
 BUF_X1 rebuffer46 (.A(\sa12_sr[0] ),
    .Z(net530));
 BUF_X4 rebuffer47 (.A(\sa12_sr[0] ),
    .Z(net531));
 BUF_X1 rebuffer48 (.A(net930),
    .Z(net532));
 BUF_X1 rebuffer49 (.A(\sa12_sr[1] ),
    .Z(net533));
 BUF_X8 rebuffer50 (.A(_04337_),
    .Z(net534));
 BUF_X8 rebuffer51 (.A(_04337_),
    .Z(net535));
 BUF_X4 rebuffer52 (.A(_14842_),
    .Z(net536));
 BUF_X1 rebuffer54 (.A(_14956_),
    .Z(net538));
 BUF_X1 rebuffer55 (.A(_06606_),
    .Z(net539));
 BUF_X4 clone56 (.A(net541),
    .Z(net540));
 BUF_X1 rebuffer57 (.A(_14993_),
    .Z(net541));
 BUF_X1 rebuffer58 (.A(_06608_),
    .Z(net542));
 BUF_X1 rebuffer59 (.A(net542),
    .Z(net543));
 BUF_X1 rebuffer60 (.A(\sa31_sub[1] ),
    .Z(net544));
 BUF_X1 rebuffer61 (.A(net595),
    .Z(net545));
 BUF_X1 rebuffer62 (.A(_12502_),
    .Z(net546));
 BUF_X1 rebuffer63 (.A(net546),
    .Z(net547));
 BUF_X1 rebuffer64 (.A(net547),
    .Z(net548));
 BUF_X1 rebuffer65 (.A(\sa12_sr[7] ),
    .Z(net549));
 BUF_X1 rebuffer66 (.A(\sa12_sr[7] ),
    .Z(net550));
 BUF_X1 rebuffer67 (.A(net550),
    .Z(net551));
 BUF_X1 rebuffer68 (.A(\sa12_sr[7] ),
    .Z(net552));
 BUF_X1 rebuffer69 (.A(_11848_),
    .Z(net553));
 BUF_X1 rebuffer70 (.A(net553),
    .Z(net554));
 BUF_X1 rebuffer71 (.A(net554),
    .Z(net555));
 BUF_X1 rebuffer72 (.A(\sa20_sub[1] ),
    .Z(net556));
 BUF_X2 rebuffer73 (.A(net556),
    .Z(net557));
 BUF_X1 rebuffer74 (.A(\sa20_sub[1] ),
    .Z(net558));
 BUF_X1 rebuffer75 (.A(\u0.tmp_w[17] ),
    .Z(net559));
 BUF_X1 rebuffer76 (.A(_03581_),
    .Z(net560));
 BUF_X1 rebuffer77 (.A(_03581_),
    .Z(net561));
 BUF_X2 split78 (.A(_14906_),
    .Z(net562));
 BUF_X1 rebuffer79 (.A(_15172_),
    .Z(net563));
 BUF_X2 rebuffer80 (.A(_15172_),
    .Z(net564));
 BUF_X1 rebuffer81 (.A(net564),
    .Z(net565));
 BUF_X8 rebuffer82 (.A(_00945_),
    .Z(net566));
 BUF_X1 rebuffer83 (.A(_09725_),
    .Z(net567));
 BUF_X1 rebuffer85 (.A(net568),
    .Z(net569));
 BUF_X1 rebuffer86 (.A(_15020_),
    .Z(net570));
 BUF_X1 rebuffer87 (.A(_15020_),
    .Z(net571));
 BUF_X1 rebuffer88 (.A(net571),
    .Z(net572));
 BUF_X1 rebuffer89 (.A(_10455_),
    .Z(net573));
 BUF_X1 rebuffer90 (.A(net573),
    .Z(net574));
 BUF_X2 rebuffer91 (.A(_14897_),
    .Z(net575));
 BUF_X1 rebuffer92 (.A(_11121_),
    .Z(net576));
 BUF_X1 rebuffer93 (.A(net576),
    .Z(net577));
 BUF_X1 rebuffer94 (.A(\sa03_sr[0] ),
    .Z(net578));
 BUF_X1 rebuffer95 (.A(\sa10_sub[0] ),
    .Z(net579));
 BUF_X1 rebuffer96 (.A(_15140_),
    .Z(net580));
 BUF_X1 rebuffer97 (.A(net580),
    .Z(net581));
 BUF_X16 clone99 (.A(net610),
    .Z(net582));
 BUF_X1 rebuffer100 (.A(\sa02_sr[1] ),
    .Z(net583));
 BUF_X1 rebuffer101 (.A(\sa02_sr[1] ),
    .Z(net584));
 BUF_X1 rebuffer102 (.A(net584),
    .Z(net585));
 BUF_X1 rebuffer103 (.A(\sa02_sr[1] ),
    .Z(net586));
 BUF_X8 clone104 (.A(_08970_),
    .Z(net587));
 BUF_X2 rebuffer105 (.A(_02389_),
    .Z(net588));
 BUF_X1 rebuffer106 (.A(_08980_),
    .Z(net589));
 BUF_X4 rebuffer108 (.A(net1192),
    .Z(net591));
 BUF_X1 rebuffer109 (.A(_01599_),
    .Z(net592));
 BUF_X1 rebuffer110 (.A(_01599_),
    .Z(net593));
 BUF_X8 clone111 (.A(_09099_),
    .Z(net594));
 BUF_X4 rebuffer112 (.A(\sa31_sub[1] ),
    .Z(net595));
 BUF_X1 rebuffer113 (.A(\sa20_sub[0] ),
    .Z(net596));
 BUF_X1 rebuffer114 (.A(\sa20_sub[0] ),
    .Z(net597));
 BUF_X4 rebuffer115 (.A(\sa20_sub[0] ),
    .Z(net598));
 BUF_X1 rebuffer117 (.A(net604),
    .Z(net600));
 BUF_X2 rebuffer613 (.A(_14706_),
    .Z(net1224));
 BUF_X1 rebuffer119 (.A(net1209),
    .Z(net602));
 BUF_X1 rebuffer120 (.A(net1209),
    .Z(net603));
 BUF_X1 rebuffer121 (.A(net1209),
    .Z(net604));
 BUF_X1 rebuffer122 (.A(net604),
    .Z(net605));
 BUF_X2 rebuffer123 (.A(_12526_),
    .Z(net606));
 BUF_X1 rebuffer124 (.A(net606),
    .Z(net607));
 BUF_X2 rebuffer125 (.A(net607),
    .Z(net608));
 BUF_X1 rebuffer126 (.A(_09153_),
    .Z(net609));
 INV_X4 clone128 (.A(net612),
    .ZN(net611));
 BUF_X4 clone129 (.A(net613),
    .Z(net612));
 BUF_X1 rebuffer130 (.A(_14989_),
    .Z(net613));
 BUF_X4 rebuffer131 (.A(_06351_),
    .Z(net614));
 BUF_X1 rebuffer133 (.A(net706),
    .Z(net616));
 BUF_X4 rebuffer135 (.A(_14838_),
    .Z(net618));
 BUF_X2 rebuffer136 (.A(_14838_),
    .Z(net619));
 BUF_X1 rebuffer137 (.A(net619),
    .Z(net620));
 BUF_X1 rebuffer152 (.A(\sa10_sr[1] ),
    .Z(net629));
 BUF_X1 rebuffer153 (.A(net629),
    .Z(net630));
 BUF_X1 rebuffer154 (.A(\sa10_sr[1] ),
    .Z(net631));
 BUF_X1 rebuffer161 (.A(\sa21_sr[1] ),
    .Z(net635));
 BUF_X1 rebuffer162 (.A(\sa21_sr[1] ),
    .Z(net636));
 BUF_X1 rebuffer163 (.A(_09717_),
    .Z(net637));
 BUF_X1 rebuffer164 (.A(net637),
    .Z(net638));
 BUF_X1 rebuffer165 (.A(_04228_),
    .Z(net639));
 BUF_X1 rebuffer166 (.A(_12623_),
    .Z(net640));
 BUF_X1 rebuffer167 (.A(\sa30_sub[0] ),
    .Z(net641));
 BUF_X1 rebuffer168 (.A(\sa30_sub[0] ),
    .Z(net642));
 BUF_X1 rebuffer169 (.A(\sa21_sr[1] ),
    .Z(net643));
 NAND3_X2 clone172 (.A1(net536),
    .A2(_09859_),
    .A3(_09861_),
    .ZN(net645));
 BUF_X4 rebuffer180 (.A(net707),
    .Z(net647));
 BUF_X4 rebuffer181 (.A(_14893_),
    .Z(net648));
 INV_X4 clone182 (.A(net650),
    .ZN(net649));
 BUF_X1 rebuffer183 (.A(net883),
    .Z(net650));
 BUF_X8 clone184 (.A(_11131_),
    .Z(net651));
 BUF_X2 clone188 (.A(net655),
    .Z(net654));
 BUF_X4 rebuffer189 (.A(_15297_),
    .Z(net655));
 BUF_X2 rebuffer190 (.A(_13842_),
    .Z(net656));
 BUF_X2 rebuffer192 (.A(\sa03_sr[1] ),
    .Z(net658));
 BUF_X4 rebuffer193 (.A(_15297_),
    .Z(net659));
 BUF_X1 rebuffer194 (.A(_11166_),
    .Z(net660));
 BUF_X1 rebuffer195 (.A(_05523_),
    .Z(net661));
 BUF_X1 rebuffer202 (.A(_14964_),
    .Z(net665));
 BUF_X1 rebuffer203 (.A(net665),
    .Z(net666));
 BUF_X1 rebuffer204 (.A(_09797_),
    .Z(net667));
 BUF_X4 rebuffer205 (.A(_09739_),
    .Z(net668));
 BUF_X2 rebuffer206 (.A(net668),
    .Z(net669));
 BUF_X1 rebuffer207 (.A(_09797_),
    .Z(net670));
 BUF_X4 rebuffer218 (.A(_15059_),
    .Z(net681));
 BUF_X2 clone219 (.A(net683),
    .Z(net682));
 BUF_X1 rebuffer220 (.A(net687),
    .Z(net683));
 BUF_X1 rebuffer221 (.A(_00939_),
    .Z(net684));
 BUF_X1 rebuffer222 (.A(_00944_),
    .Z(net685));
 BUF_X2 rebuffer223 (.A(_01241_),
    .Z(net686));
 BUF_X4 rebuffer224 (.A(_15053_),
    .Z(net687));
 BUF_X1 rebuffer226 (.A(_09733_),
    .Z(net689));
 BUF_X4 rebuffer227 (.A(_03585_),
    .Z(net690));
 BUF_X1 rebuffer228 (.A(_11856_),
    .Z(net691));
 BUF_X2 rebuffer229 (.A(_11856_),
    .Z(net692));
 BUF_X8 rebuffer230 (.A(_03672_),
    .Z(net693));
 BUF_X1 rebuffer231 (.A(\sa20_sr[1] ),
    .Z(net694));
 BUF_X1 rebuffer232 (.A(net694),
    .Z(net695));
 BUF_X1 rebuffer233 (.A(net694),
    .Z(net696));
 BUF_X4 rebuffer245 (.A(_05177_),
    .Z(net708));
 BUF_X1 rebuffer246 (.A(_15274_),
    .Z(net709));
 BUF_X1 rebuffer247 (.A(_13224_),
    .Z(net710));
 BUF_X1 rebuffer248 (.A(_10437_),
    .Z(net711));
 BUF_X4 rebuffer249 (.A(_10506_),
    .Z(net712));
 BUF_X4 clone257 (.A(net721),
    .Z(net720));
 BUF_X1 rebuffer258 (.A(net730),
    .Z(net721));
 INV_X4 clone259 (.A(_12506_),
    .ZN(net722));
 BUF_X8 clone260 (.A(_12508_),
    .Z(net723));
 BUF_X4 clone262 (.A(net726),
    .Z(net725));
 BUF_X2 rebuffer263 (.A(_15161_),
    .Z(net726));
 BUF_X4 clone264 (.A(_02936_),
    .Z(net727));
 BUF_X4 clone271 (.A(net10),
    .Z(net734));
 BUF_X4 rebuffer274 (.A(_01086_),
    .Z(net737));
 BUF_X8 rebuffer275 (.A(_01227_),
    .Z(net738));
 BUF_X1 rebuffer276 (.A(net738),
    .Z(net739));
 BUF_X4 clone277 (.A(net1030),
    .Z(net740));
 BUF_X8 clone278 (.A(_00946_),
    .Z(net741));
 BUF_X8 clone279 (.A(net844),
    .Z(net742));
 BUF_X8 rebuffer280 (.A(_01086_),
    .Z(net743));
 BUF_X2 rebuffer281 (.A(_15210_),
    .Z(net744));
 BUF_X4 rebuffer282 (.A(_15196_),
    .Z(net745));
 BUF_X1 rebuffer283 (.A(net745),
    .Z(net746));
 BUF_X1 rebuffer284 (.A(_03580_),
    .Z(net747));
 BUF_X1 rebuffer289 (.A(\sa01_sr[1] ),
    .Z(net752));
 BUF_X1 rebuffer290 (.A(\sa01_sr[1] ),
    .Z(net753));
 BUF_X1 rebuffer291 (.A(\sa30_sub[1] ),
    .Z(net754));
 BUF_X1 rebuffer292 (.A(\sa30_sub[1] ),
    .Z(net755));
 BUF_X4 rebuffer293 (.A(_15095_),
    .Z(net756));
 BUF_X4 rebuffer294 (.A(_01708_),
    .Z(net757));
 BUF_X2 rebuffer295 (.A(net757),
    .Z(net758));
 BUF_X4 rebuffer296 (.A(\sa21_sr[0] ),
    .Z(net759));
 BUF_X1 rebuffer297 (.A(net759),
    .Z(net760));
 BUF_X4 clone298 (.A(net762),
    .Z(net761));
 BUF_X1 rebuffer299 (.A(_15095_),
    .Z(net762));
 BUF_X8 clone300 (.A(_01604_),
    .Z(net763));
 BUF_X4 rebuffer301 (.A(_04479_),
    .Z(net764));
 BUF_X1 rebuffer302 (.A(_04232_),
    .Z(net765));
 BUF_X1 rebuffer303 (.A(net765),
    .Z(net766));
 BUF_X1 rebuffer304 (.A(net765),
    .Z(net767));
 BUF_X4 rebuffer305 (.A(net777),
    .Z(net768));
 BUF_X2 rebuffer306 (.A(net777),
    .Z(net769));
 BUF_X1 rebuffer307 (.A(net777),
    .Z(net770));
 BUF_X1 rebuffer308 (.A(net1202),
    .Z(net771));
 BUF_X4 rebuffer309 (.A(_04233_),
    .Z(net772));
 BUF_X1 rebuffer310 (.A(net772),
    .Z(net773));
 BUF_X1 rebuffer311 (.A(_09717_),
    .Z(net774));
 BUF_X1 split312 (.A(_15242_),
    .Z(net775));
 BUF_X16 clone313 (.A(_04388_),
    .Z(net776));
 BUF_X4 rebuffer314 (.A(_15230_),
    .Z(net777));
 BUF_X1 rebuffer315 (.A(net777),
    .Z(net778));
 BUF_X2 rebuffer316 (.A(_04351_),
    .Z(net779));
 BUF_X1 rebuffer317 (.A(_04351_),
    .Z(net780));
 BUF_X1 rebuffer320 (.A(net782),
    .Z(net783));
 BUF_X1 rebuffer321 (.A(net782),
    .Z(net784));
 BUF_X1 rebuffer322 (.A(\u0.w[1][24] ),
    .Z(net785));
 BUF_X1 rebuffer324 (.A(\u0.tmp_w[24] ),
    .Z(net787));
 BUF_X1 rebuffer325 (.A(\u0.tmp_w[24] ),
    .Z(net788));
 BUF_X8 rebuffer326 (.A(_14776_),
    .Z(net789));
 BUF_X1 rebuffer327 (.A(_06625_),
    .Z(net790));
 BUF_X4 rebuffer328 (.A(net1234),
    .Z(net791));
 BUF_X2 rebuffer329 (.A(net791),
    .Z(net792));
 BUF_X1 rebuffer330 (.A(_06604_),
    .Z(net793));
 BUF_X1 rebuffer331 (.A(net793),
    .Z(net794));
 BUF_X1 rebuffer333 (.A(\u0.w[2][25] ),
    .Z(net796));
 BUF_X2 rebuffer334 (.A(net796),
    .Z(net797));
 BUF_X1 rebuffer335 (.A(net797),
    .Z(net798));
 BUF_X1 rebuffer353 (.A(_05013_),
    .Z(net816));
 BUF_X8 rebuffer354 (.A(_15265_),
    .Z(net817));
 BUF_X2 rebuffer355 (.A(net817),
    .Z(net818));
 BUF_X1 rebuffer356 (.A(net817),
    .Z(net819));
 BUF_X4 rebuffer362 (.A(net826),
    .Z(net825));
 BUF_X4 rebuffer363 (.A(_14810_),
    .Z(net826));
 BUF_X8 rebuffer364 (.A(_09129_),
    .Z(net827));
 BUF_X2 rebuffer367 (.A(_15242_),
    .Z(net830));
 BUF_X1 rebuffer374 (.A(\sa00_sr[1] ),
    .Z(net837));
 BUF_X1 rebuffer375 (.A(net837),
    .Z(net838));
 BUF_X1 rebuffer376 (.A(\sa00_sr[1] ),
    .Z(net839));
 BUF_X1 rebuffer377 (.A(_11843_),
    .Z(net840));
 BUF_X8 rebuffer378 (.A(_11852_),
    .Z(net841));
 BUF_X1 rebuffer379 (.A(net841),
    .Z(net842));
 BUF_X1 rebuffer385 (.A(_14874_),
    .Z(net848));
 BUF_X1 rebuffer408 (.A(net870),
    .Z(net871));
 BUF_X1 rebuffer422 (.A(net884),
    .Z(net885));
 BUF_X4 rebuffer433 (.A(_15262_),
    .Z(net896));
 BUF_X1 rebuffer434 (.A(net896),
    .Z(net897));
 BUF_X1 rebuffer435 (.A(_15270_),
    .Z(net898));
 BUF_X8 clone438 (.A(net836),
    .Z(net901));
 BUF_X4 clone439 (.A(_05663_),
    .Z(net902));
 BUF_X4 rebuffer446 (.A(_15306_),
    .Z(net909));
 BUF_X8 clone447 (.A(_05548_),
    .Z(net910));
 BUF_X4 rebuffer456 (.A(\sa30_sr[0] ),
    .Z(net919));
 BUF_X1 rebuffer457 (.A(\sa30_sr[0] ),
    .Z(net920));
 BUF_X1 rebuffer458 (.A(\sa30_sr[0] ),
    .Z(net921));
 BUF_X1 rebuffer459 (.A(_08983_),
    .Z(net922));
 BUF_X4 rebuffer460 (.A(_15057_),
    .Z(net923));
 BUF_X1 rebuffer461 (.A(net923),
    .Z(net924));
 BUF_X4 clone462 (.A(net926),
    .Z(net925));
 BUF_X1 rebuffer463 (.A(_15054_),
    .Z(net926));
 BUF_X4 rebuffer468 (.A(_14970_),
    .Z(net931));
 BUF_X1 rebuffer469 (.A(net931),
    .Z(net932));
 BUF_X1 rebuffer480 (.A(_15206_),
    .Z(net943));
 BUF_X1 rebuffer481 (.A(net943),
    .Z(net944));
 BUF_X1 rebuffer496 (.A(_11123_),
    .Z(net959));
 BUF_X4 clone497 (.A(net961),
    .Z(net960));
 BUF_X1 rebuffer498 (.A(_13839_),
    .Z(net961));
 BUF_X2 rebuffer499 (.A(_13875_),
    .Z(net962));
 BUF_X1 rebuffer500 (.A(net962),
    .Z(net963));
 BUF_X1 rebuffer501 (.A(_13875_),
    .Z(net964));
 BUF_X1 rebuffer502 (.A(_13875_),
    .Z(net965));
 BUF_X1 rebuffer503 (.A(_11137_),
    .Z(net966));
 BUF_X4 rebuffer504 (.A(_15025_),
    .Z(net967));
 BUF_X4 rebuffer505 (.A(_15025_),
    .Z(net968));
 BUF_X8 rebuffer506 (.A(_13926_),
    .Z(net969));
 BUF_X1 rebuffer507 (.A(_13832_),
    .Z(net970));
 BUF_X1 rebuffer508 (.A(\sa32_sub[1] ),
    .Z(net971));
 BUF_X1 rebuffer509 (.A(_11122_),
    .Z(net972));
 BUF_X1 rebuffer510 (.A(net972),
    .Z(net973));
 BUF_X2 rebuffer511 (.A(\sa32_sub[1] ),
    .Z(net974));
 BUF_X2 rebuffer514 (.A(net979),
    .Z(net977));
 BUF_X4 clone515 (.A(net980),
    .Z(net978));
 BUF_X4 rebuffer516 (.A(_14929_),
    .Z(net979));
 BUF_X1 rebuffer517 (.A(_14929_),
    .Z(net980));
 BUF_X1 rebuffer518 (.A(_11946_),
    .Z(net981));
 BUF_X2 rebuffer522 (.A(_14865_),
    .Z(net985));
 BUF_X1 rebuffer523 (.A(_10802_),
    .Z(net986));
 BUF_X4 clone524 (.A(net988),
    .Z(net987));
 BUF_X1 rebuffer525 (.A(net989),
    .Z(net988));
 BUF_X1 rebuffer526 (.A(_10450_),
    .Z(net989));
 BUF_X4 rebuffer538 (.A(_14772_),
    .Z(net1001));
 BUF_X1 rebuffer539 (.A(_14772_),
    .Z(net1002));
 BUF_X1 rebuffer548 (.A(_12114_),
    .Z(net1011));
 AOI21_X2 clone549 (.A(_11969_),
    .B1(_11925_),
    .B2(_11930_),
    .ZN(net1012));
 BUF_X8 clone550 (.A(_12052_),
    .Z(net1013));
 BUF_X16 clone551 (.A(net715),
    .Z(net1014));
 BUF_X1 rebuffer553 (.A(_06334_),
    .Z(net1016));
 BUF_X1 rebuffer554 (.A(\u0.tmp_w[1] ),
    .Z(net1017));
 BUF_X1 rebuffer555 (.A(net1017),
    .Z(net1018));
 BUF_X1 rebuffer556 (.A(\u0.tmp_w[0] ),
    .Z(net1019));
 BUF_X1 rebuffer557 (.A(net1019),
    .Z(net1020));
 BUF_X1 rebuffer558 (.A(net1019),
    .Z(net1021));
 BUF_X4 rebuffer570 (.A(_15066_),
    .Z(net1033));
 BUF_X8 rebuffer573 (.A(_03777_),
    .Z(net1036));
 BUF_X4 rebuffer576 (.A(_02463_),
    .Z(net1039));
 BUF_X4 clone577 (.A(_02279_),
    .Z(net1040));
 BUF_X16 rebuffer578 (.A(net729),
    .Z(net1041));
 BUF_X8 rebuffer579 (.A(_15140_),
    .Z(net1042));
 BUF_X1 rebuffer580 (.A(net1042),
    .Z(net1043));
 BUF_X8 clone581 (.A(net731),
    .Z(net1044));
 BUF_X1 rebuffer586 (.A(\u0.tmp_w[9] ),
    .Z(net1049));
 BUF_X1 rebuffer587 (.A(\u0.subword[9] ),
    .Z(net1050));
 BUF_X8 rebuffer588 (.A(_07434_),
    .Z(net1051));
 BUF_X2 rebuffer589 (.A(net1051),
    .Z(net1052));
 BUF_X2 rebuffer590 (.A(net1051),
    .Z(net1053));
 BUF_X1 rebuffer591 (.A(net1227),
    .Z(net1054));
 BUF_X4 clone593 (.A(net1057),
    .Z(net1056));
 BUF_X1 rebuffer594 (.A(net942),
    .Z(net1057));
 BUF_X1 rebuffer605 (.A(\sa31_sub[1] ),
    .Z(net1068));
 BUF_X1 rebuffer606 (.A(\sa12_sr[0] ),
    .Z(net1069));
 BUF_X4 rebuffer614 (.A(_04265_),
    .Z(net1077));
 BUF_X1 rebuffer615 (.A(net1077),
    .Z(net1078));
 BUF_X1 rebuffer616 (.A(net1077),
    .Z(net1079));
 BUF_X1 rebuffer617 (.A(net1077),
    .Z(net1080));
 BUF_X1 rebuffer618 (.A(net1080),
    .Z(net1081));
 BUF_X1 rebuffer619 (.A(_04265_),
    .Z(net1082));
 BUF_X1 rebuffer625 (.A(net1087),
    .Z(net1088));
 BUF_X1 rebuffer626 (.A(net1087),
    .Z(net1089));
 BUF_X1 rebuffer632 (.A(_02310_),
    .Z(net1095));
 BUF_X1 rebuffer633 (.A(net1095),
    .Z(net1096));
 BUF_X4 rebuffer634 (.A(_02643_),
    .Z(net1097));
 BUF_X2 rebuffer636 (.A(_12017_),
    .Z(net1099));
 BUF_X1 rebuffer637 (.A(net1099),
    .Z(net1100));
 BUF_X1 rebuffer638 (.A(_11843_),
    .Z(net1101));
 BUF_X1 rebuffer639 (.A(_09006_),
    .Z(net1102));
 BUF_X1 rebuffer640 (.A(net1102),
    .Z(net1103));
 BUF_X2 rebuffer641 (.A(_09006_),
    .Z(net1104));
 OAI21_X2 clone649 (.A(_05092_),
    .B1(_04940_),
    .B2(_04946_),
    .ZN(net1112));
 BUF_X2 rebuffer651 (.A(_15265_),
    .Z(net1114));
 BUF_X2 rebuffer654 (.A(net1169),
    .Z(net1117));
 BUF_X2 rebuffer655 (.A(_14730_),
    .Z(net1118));
 BUF_X2 rebuffer656 (.A(net1118),
    .Z(net1119));
 BUF_X1 rebuffer657 (.A(net1119),
    .Z(net1120));
 BUF_X1 rebuffer658 (.A(net1119),
    .Z(net1121));
 BUF_X4 rebuffer659 (.A(net1182),
    .Z(net1122));
 BUF_X1 rebuffer660 (.A(net1122),
    .Z(net1123));
 BUF_X4 rebuffer667 (.A(_01862_),
    .Z(net1130));
 BUF_X2 rebuffer668 (.A(net1130),
    .Z(net1131));
 BUF_X4 rebuffer669 (.A(net1130),
    .Z(net1132));
 BUF_X2 clone670 (.A(net1134),
    .Z(net1133));
 BUF_X1 rebuffer671 (.A(_15098_),
    .Z(net1134));
 BUF_X1 rebuffer685 (.A(_04897_),
    .Z(net1148));
 BUF_X1 rebuffer686 (.A(_04928_),
    .Z(net1149));
 BUF_X1 rebuffer687 (.A(_04928_),
    .Z(net1150));
 BUF_X1 rebuffer688 (.A(net1150),
    .Z(net1151));
 BUF_X1 rebuffer689 (.A(net1151),
    .Z(net1152));
 BUF_X8 clone690 (.A(net1154),
    .Z(net1153));
 BUF_X1 rebuffer691 (.A(_04863_),
    .Z(net1154));
 BUF_X4 clone692 (.A(net1156),
    .Z(net1155));
 BUF_X2 clone693 (.A(_15261_),
    .Z(net1156));
 INV_X4 clone694 (.A(net698),
    .ZN(net1157));
 BUF_X1 rebuffer695 (.A(_04863_),
    .Z(net1158));
 BUF_X4 clone700 (.A(net1164),
    .Z(net1163));
 BUF_X1 rebuffer701 (.A(_14735_),
    .Z(net1164));
 BUF_X1 rebuffer704 (.A(net1166),
    .Z(net1167));
 BUF_X1 rebuffer711 (.A(_02348_),
    .Z(net1174));
 BUF_X2 rebuffer712 (.A(net1174),
    .Z(net1175));
 BUF_X4 clone720 (.A(net1184),
    .Z(net1183));
 BUF_X1 rebuffer721 (.A(_15034_),
    .Z(net1184));
 BUF_X4 clone722 (.A(_13840_),
    .Z(net1185));
 BUF_X4 rebuffer723 (.A(_13839_),
    .Z(net1186));
 BUF_X8 clone724 (.A(_13840_),
    .Z(net1187));
 BUF_X1 rebuffer725 (.A(_13941_),
    .Z(net1188));
 BUF_X1 rebuffer731 (.A(_14665_),
    .Z(net1194));
 BUF_X1 rebuffer732 (.A(_14676_),
    .Z(net1195));
 BUF_X1 rebuffer733 (.A(net1195),
    .Z(net1196));
 BUF_X2 rebuffer737 (.A(_14926_),
    .Z(net1200));
 BUF_X4 rebuffer738 (.A(_15104_),
    .Z(net1201));
 BUF_X8 clone742 (.A(_06868_),
    .Z(net1205));
 BUF_X2 rebuffer743 (.A(_13996_),
    .Z(net1206));
 BUF_X1 rebuffer744 (.A(_15022_),
    .Z(net1207));
 BUF_X1 rebuffer768 (.A(_14694_),
    .Z(net1231));
 INV_X4 clone769 (.A(_07426_),
    .ZN(net1232));
 BUF_X4 rebuffer770 (.A(_06475_),
    .Z(net1233));
 BUF_X1 rebuffer773 (.A(_06460_),
    .Z(net1236));
 BUF_X1 rebuffer774 (.A(_07448_),
    .Z(net1237));
 BUF_X2 split775 (.A(_14701_),
    .Z(net1238));
 BUF_X1 rebuffer56 (.A(_13284_),
    .Z(net1));
 BUF_X1 rebuffer78 (.A(_06265_),
    .Z(net615));
 BUF_X1 rebuffer98 (.A(\sa20_sub[0] ),
    .Z(net621));
 BUF_X2 rebuffer159 (.A(_12732_),
    .Z(net673));
 BUF_X8 rebuffer188 (.A(_04972_),
    .Z(net698));
 BUF_X4 rebuffer208 (.A(\sa11_sr[7] ),
    .Z(net705));
 BUF_X1 rebuffer209 (.A(net705),
    .Z(net706));
 BUF_X4 rebuffer210 (.A(_14833_),
    .Z(net707));
 BUF_X1 rebuffer212 (.A(_11844_),
    .Z(net714));
 BUF_X1 rebuffer216 (.A(_15131_),
    .Z(net718));
 BUF_X2 rebuffer217 (.A(_02423_),
    .Z(net719));
 BUF_X4 rebuffer225 (.A(_02341_),
    .Z(net728));
 BUF_X4 rebuffer234 (.A(_02278_),
    .Z(net729));
 BUF_X1 rebuffer235 (.A(net729),
    .Z(net730));
 INV_X4 clone236 (.A(net1041),
    .ZN(net731));
 BUF_X4 clone237 (.A(net735),
    .Z(net732));
 BUF_X1 rebuffer238 (.A(_15129_),
    .Z(net735));
 BUF_X1 rebuffer250 (.A(_06252_),
    .Z(net802));
 BUF_X1 rebuffer251 (.A(_04479_),
    .Z(net803));
 BUF_X1 rebuffer253 (.A(_01872_),
    .Z(net805));
 BUF_X2 rebuffer255 (.A(_01706_),
    .Z(net807));
 BUF_X1 rebuffer277 (.A(_07902_),
    .Z(net829));
 BUF_X8 clone280 (.A(net827),
    .Z(net831));
 BUF_X16 clone281 (.A(_09209_),
    .Z(net832));
 BUF_X8 rebuffer287 (.A(_00945_),
    .Z(net835));
 INV_X4 clone299 (.A(net835),
    .ZN(net844));
 BUF_X4 rebuffer312 (.A(_15201_),
    .Z(net847));
 BUF_X8 clone314 (.A(_03586_),
    .Z(net850));
 BUF_X1 rebuffer318 (.A(_14897_),
    .Z(net851));
 BUF_X2 rebuffer336 (.A(_14897_),
    .Z(net852));
 BUF_X1 rebuffer365 (.A(_14828_),
    .Z(net879));
 BUF_X2 rebuffer395 (.A(_12683_),
    .Z(net911));
 BUF_X1 rebuffer399 (.A(net914),
    .Z(net915));
 BUF_X8 clone400 (.A(_04234_),
    .Z(net916));
 BUF_X1 rebuffer402 (.A(_12209_),
    .Z(net918));
 BUF_X4 clone408 (.A(net935),
    .Z(net934));
 BUF_X1 rebuffer409 (.A(_09733_),
    .Z(net935));
 BUF_X4 rebuffer410 (.A(_09733_),
    .Z(net936));
 BUF_X8 rebuffer411 (.A(_00977_),
    .Z(net937));
 BUF_X1 rebuffer412 (.A(net937),
    .Z(net938));
 BUF_X1 rebuffer413 (.A(net937),
    .Z(net939));
 BUF_X4 rebuffer414 (.A(net937),
    .Z(net940));
 BUF_X4 rebuffer415 (.A(_00960_),
    .Z(net941));
 BUF_X2 rebuffer416 (.A(_15064_),
    .Z(net942));
 BUF_X1 rebuffer418 (.A(_09153_),
    .Z(net946));
 BUF_X16 clone419 (.A(_09010_),
    .Z(net947));
 BUF_X16 clone420 (.A(_09009_),
    .Z(net948));
 BUF_X16 clone421 (.A(_09011_),
    .Z(net949));
 BUF_X16 clone422 (.A(_00962_),
    .Z(net950));
 BUF_X16 clone423 (.A(_09012_),
    .Z(net951));
 BUF_X2 rebuffer427 (.A(_14708_),
    .Z(net955));
 BUF_X1 rebuffer428 (.A(net955),
    .Z(net956));
 BUF_X8 clone437 (.A(net993),
    .Z(net992));
 BUF_X1 rebuffer438 (.A(_06609_),
    .Z(net993));
 BUF_X4 rebuffer443 (.A(_09979_),
    .Z(net997));
 BUF_X8 clone445 (.A(_06319_),
    .Z(net999));
 BUF_X4 clone446 (.A(_06253_),
    .Z(net1000));
 BUF_X4 clone448 (.A(net1004),
    .Z(net1003));
 BUF_X1 rebuffer449 (.A(\u0.w[0][18] ),
    .Z(net1004));
 INV_X4 clone472 (.A(net835),
    .ZN(net1030));
 BUF_X8 rebuffer476 (.A(_02967_),
    .Z(net1037));
 BUF_X1 rebuffer477 (.A(net1037),
    .Z(net1038));
 BUF_X4 clone478 (.A(net1046),
    .Z(net1045));
 BUF_X1 rebuffer479 (.A(_15162_),
    .Z(net1046));
 BUF_X8 clone514 (.A(_02953_),
    .Z(net1084));
 BUF_X16 clone516 (.A(_09099_),
    .Z(net1085));
 BUF_X16 clone532 (.A(_06611_),
    .Z(net1116));
 INV_X16 clone533 (.A(_06610_),
    .ZN(net1124));
 INV_X4 clone547 (.A(net841),
    .ZN(net1144));
 BUF_X1 rebuffer559 (.A(_14796_),
    .Z(net1147));
 BUF_X1 rebuffer560 (.A(_14796_),
    .Z(net1159));
 BUF_X1 rebuffer564 (.A(_06355_),
    .Z(net1165));
 BUF_X4 clone565 (.A(_06378_),
    .Z(net1168));
 BUF_X4 rebuffer566 (.A(_14730_),
    .Z(net1169));
 BUF_X1 rebuffer567 (.A(net1169),
    .Z(net1170));
 BUF_X1 rebuffer581 (.A(_14733_),
    .Z(net1182));
 BUF_X4 rebuffer582 (.A(_04567_),
    .Z(net1189));
 BUF_X2 rebuffer583 (.A(_04567_),
    .Z(net1190));
 BUF_X2 rebuffer584 (.A(net1190),
    .Z(net1191));
 BUF_X4 rebuffer592 (.A(_15233_),
    .Z(net1192));
 BUF_X1 rebuffer593 (.A(_15233_),
    .Z(net1197));
 BUF_X1 rebuffer595 (.A(net1197),
    .Z(net1198));
 BUF_X2 rebuffer596 (.A(_15230_),
    .Z(net1202));
 BUF_X16 clone597 (.A(_04235_),
    .Z(net1203));
 BUF_X4 rebuffer599 (.A(_06335_),
    .Z(net1209));
 BUF_X1 rebuffer621 (.A(net1225),
    .Z(net1226));
 BUF_X1 rebuffer622 (.A(_06460_),
    .Z(net1227));
 BUF_X4 rebuffer628 (.A(_14767_),
    .Z(net1230));
 BUF_X2 rebuffer629 (.A(_14767_),
    .Z(net1234));
 BUF_X16 clone630 (.A(_06612_),
    .Z(net1235));
 INV_X2 clone631 (.A(net1241),
    .ZN(net1240));
 BUF_X1 rebuffer642 (.A(_14701_),
    .Z(net1241));
 FILLCELL_X32 FILLER_0_1 ();
 FILLCELL_X32 FILLER_0_33 ();
 FILLCELL_X32 FILLER_0_65 ();
 FILLCELL_X32 FILLER_0_97 ();
 FILLCELL_X32 FILLER_0_129 ();
 FILLCELL_X32 FILLER_0_161 ();
 FILLCELL_X32 FILLER_0_193 ();
 FILLCELL_X32 FILLER_0_225 ();
 FILLCELL_X32 FILLER_0_257 ();
 FILLCELL_X32 FILLER_0_289 ();
 FILLCELL_X32 FILLER_0_321 ();
 FILLCELL_X16 FILLER_0_353 ();
 FILLCELL_X32 FILLER_0_374 ();
 FILLCELL_X32 FILLER_0_406 ();
 FILLCELL_X16 FILLER_0_438 ();
 FILLCELL_X2 FILLER_0_454 ();
 FILLCELL_X4 FILLER_0_463 ();
 FILLCELL_X2 FILLER_0_467 ();
 FILLCELL_X2 FILLER_0_473 ();
 FILLCELL_X1 FILLER_0_475 ();
 FILLCELL_X2 FILLER_0_489 ();
 FILLCELL_X2 FILLER_0_514 ();
 FILLCELL_X1 FILLER_0_516 ();
 FILLCELL_X1 FILLER_0_532 ();
 FILLCELL_X2 FILLER_0_536 ();
 FILLCELL_X1 FILLER_0_538 ();
 FILLCELL_X2 FILLER_0_542 ();
 FILLCELL_X1 FILLER_0_544 ();
 FILLCELL_X2 FILLER_0_554 ();
 FILLCELL_X1 FILLER_0_556 ();
 FILLCELL_X1 FILLER_0_602 ();
 FILLCELL_X4 FILLER_0_654 ();
 FILLCELL_X1 FILLER_0_658 ();
 FILLCELL_X2 FILLER_0_662 ();
 FILLCELL_X1 FILLER_0_664 ();
 FILLCELL_X1 FILLER_0_674 ();
 FILLCELL_X1 FILLER_0_679 ();
 FILLCELL_X4 FILLER_0_703 ();
 FILLCELL_X1 FILLER_0_707 ();
 FILLCELL_X8 FILLER_0_711 ();
 FILLCELL_X1 FILLER_0_719 ();
 FILLCELL_X16 FILLER_0_724 ();
 FILLCELL_X2 FILLER_0_740 ();
 FILLCELL_X1 FILLER_0_742 ();
 FILLCELL_X8 FILLER_0_746 ();
 FILLCELL_X32 FILLER_0_761 ();
 FILLCELL_X32 FILLER_0_793 ();
 FILLCELL_X16 FILLER_0_825 ();
 FILLCELL_X8 FILLER_0_841 ();
 FILLCELL_X2 FILLER_0_849 ();
 FILLCELL_X16 FILLER_0_868 ();
 FILLCELL_X4 FILLER_0_884 ();
 FILLCELL_X1 FILLER_0_888 ();
 FILLCELL_X1 FILLER_0_905 ();
 FILLCELL_X2 FILLER_0_909 ();
 FILLCELL_X1 FILLER_0_921 ();
 FILLCELL_X16 FILLER_0_926 ();
 FILLCELL_X8 FILLER_0_942 ();
 FILLCELL_X16 FILLER_0_957 ();
 FILLCELL_X2 FILLER_0_973 ();
 FILLCELL_X4 FILLER_0_985 ();
 FILLCELL_X2 FILLER_0_989 ();
 FILLCELL_X32 FILLER_0_994 ();
 FILLCELL_X32 FILLER_0_1026 ();
 FILLCELL_X32 FILLER_0_1058 ();
 FILLCELL_X32 FILLER_0_1090 ();
 FILLCELL_X32 FILLER_0_1122 ();
 FILLCELL_X32 FILLER_0_1154 ();
 FILLCELL_X16 FILLER_0_1186 ();
 FILLCELL_X4 FILLER_0_1202 ();
 FILLCELL_X2 FILLER_0_1206 ();
 FILLCELL_X1 FILLER_0_1208 ();
 FILLCELL_X32 FILLER_1_1 ();
 FILLCELL_X32 FILLER_1_33 ();
 FILLCELL_X32 FILLER_1_65 ();
 FILLCELL_X32 FILLER_1_97 ();
 FILLCELL_X32 FILLER_1_129 ();
 FILLCELL_X32 FILLER_1_161 ();
 FILLCELL_X32 FILLER_1_193 ();
 FILLCELL_X32 FILLER_1_225 ();
 FILLCELL_X32 FILLER_1_257 ();
 FILLCELL_X32 FILLER_1_289 ();
 FILLCELL_X32 FILLER_1_321 ();
 FILLCELL_X32 FILLER_1_353 ();
 FILLCELL_X32 FILLER_1_385 ();
 FILLCELL_X32 FILLER_1_417 ();
 FILLCELL_X8 FILLER_1_449 ();
 FILLCELL_X2 FILLER_1_457 ();
 FILLCELL_X32 FILLER_1_462 ();
 FILLCELL_X16 FILLER_1_494 ();
 FILLCELL_X4 FILLER_1_510 ();
 FILLCELL_X2 FILLER_1_514 ();
 FILLCELL_X1 FILLER_1_516 ();
 FILLCELL_X4 FILLER_1_523 ();
 FILLCELL_X1 FILLER_1_527 ();
 FILLCELL_X8 FILLER_1_537 ();
 FILLCELL_X2 FILLER_1_545 ();
 FILLCELL_X1 FILLER_1_547 ();
 FILLCELL_X2 FILLER_1_551 ();
 FILLCELL_X4 FILLER_1_556 ();
 FILLCELL_X1 FILLER_1_560 ();
 FILLCELL_X1 FILLER_1_578 ();
 FILLCELL_X4 FILLER_1_583 ();
 FILLCELL_X16 FILLER_1_591 ();
 FILLCELL_X2 FILLER_1_607 ();
 FILLCELL_X2 FILLER_1_612 ();
 FILLCELL_X2 FILLER_1_617 ();
 FILLCELL_X2 FILLER_1_629 ();
 FILLCELL_X2 FILLER_1_653 ();
 FILLCELL_X8 FILLER_1_659 ();
 FILLCELL_X1 FILLER_1_667 ();
 FILLCELL_X4 FILLER_1_686 ();
 FILLCELL_X2 FILLER_1_700 ();
 FILLCELL_X1 FILLER_1_702 ();
 FILLCELL_X2 FILLER_1_729 ();
 FILLCELL_X1 FILLER_1_731 ();
 FILLCELL_X32 FILLER_1_735 ();
 FILLCELL_X32 FILLER_1_767 ();
 FILLCELL_X32 FILLER_1_799 ();
 FILLCELL_X32 FILLER_1_831 ();
 FILLCELL_X8 FILLER_1_863 ();
 FILLCELL_X2 FILLER_1_871 ();
 FILLCELL_X1 FILLER_1_873 ();
 FILLCELL_X2 FILLER_1_888 ();
 FILLCELL_X2 FILLER_1_909 ();
 FILLCELL_X4 FILLER_1_916 ();
 FILLCELL_X2 FILLER_1_920 ();
 FILLCELL_X4 FILLER_1_926 ();
 FILLCELL_X1 FILLER_1_930 ();
 FILLCELL_X2 FILLER_1_967 ();
 FILLCELL_X1 FILLER_1_969 ();
 FILLCELL_X2 FILLER_1_988 ();
 FILLCELL_X1 FILLER_1_990 ();
 FILLCELL_X4 FILLER_1_996 ();
 FILLCELL_X32 FILLER_1_1020 ();
 FILLCELL_X32 FILLER_1_1052 ();
 FILLCELL_X32 FILLER_1_1084 ();
 FILLCELL_X32 FILLER_1_1116 ();
 FILLCELL_X32 FILLER_1_1148 ();
 FILLCELL_X16 FILLER_1_1180 ();
 FILLCELL_X8 FILLER_1_1196 ();
 FILLCELL_X4 FILLER_1_1204 ();
 FILLCELL_X1 FILLER_1_1208 ();
 FILLCELL_X32 FILLER_2_1 ();
 FILLCELL_X32 FILLER_2_33 ();
 FILLCELL_X32 FILLER_2_65 ();
 FILLCELL_X32 FILLER_2_97 ();
 FILLCELL_X32 FILLER_2_129 ();
 FILLCELL_X32 FILLER_2_161 ();
 FILLCELL_X32 FILLER_2_193 ();
 FILLCELL_X32 FILLER_2_225 ();
 FILLCELL_X32 FILLER_2_257 ();
 FILLCELL_X32 FILLER_2_289 ();
 FILLCELL_X32 FILLER_2_321 ();
 FILLCELL_X32 FILLER_2_353 ();
 FILLCELL_X32 FILLER_2_385 ();
 FILLCELL_X32 FILLER_2_417 ();
 FILLCELL_X32 FILLER_2_449 ();
 FILLCELL_X32 FILLER_2_481 ();
 FILLCELL_X8 FILLER_2_513 ();
 FILLCELL_X2 FILLER_2_521 ();
 FILLCELL_X1 FILLER_2_523 ();
 FILLCELL_X16 FILLER_2_527 ();
 FILLCELL_X4 FILLER_2_543 ();
 FILLCELL_X2 FILLER_2_547 ();
 FILLCELL_X1 FILLER_2_549 ();
 FILLCELL_X16 FILLER_2_553 ();
 FILLCELL_X2 FILLER_2_569 ();
 FILLCELL_X1 FILLER_2_571 ();
 FILLCELL_X32 FILLER_2_575 ();
 FILLCELL_X2 FILLER_2_607 ();
 FILLCELL_X1 FILLER_2_632 ();
 FILLCELL_X8 FILLER_2_650 ();
 FILLCELL_X1 FILLER_2_658 ();
 FILLCELL_X32 FILLER_2_713 ();
 FILLCELL_X32 FILLER_2_745 ();
 FILLCELL_X32 FILLER_2_777 ();
 FILLCELL_X32 FILLER_2_809 ();
 FILLCELL_X16 FILLER_2_841 ();
 FILLCELL_X8 FILLER_2_857 ();
 FILLCELL_X4 FILLER_2_865 ();
 FILLCELL_X2 FILLER_2_869 ();
 FILLCELL_X4 FILLER_2_878 ();
 FILLCELL_X1 FILLER_2_882 ();
 FILLCELL_X4 FILLER_2_897 ();
 FILLCELL_X1 FILLER_2_901 ();
 FILLCELL_X2 FILLER_2_905 ();
 FILLCELL_X1 FILLER_2_907 ();
 FILLCELL_X4 FILLER_2_917 ();
 FILLCELL_X1 FILLER_2_921 ();
 FILLCELL_X4 FILLER_2_936 ();
 FILLCELL_X4 FILLER_2_969 ();
 FILLCELL_X1 FILLER_2_973 ();
 FILLCELL_X2 FILLER_2_993 ();
 FILLCELL_X4 FILLER_2_999 ();
 FILLCELL_X2 FILLER_2_1003 ();
 FILLCELL_X1 FILLER_2_1024 ();
 FILLCELL_X32 FILLER_2_1035 ();
 FILLCELL_X32 FILLER_2_1067 ();
 FILLCELL_X32 FILLER_2_1099 ();
 FILLCELL_X32 FILLER_2_1131 ();
 FILLCELL_X32 FILLER_2_1163 ();
 FILLCELL_X8 FILLER_2_1195 ();
 FILLCELL_X4 FILLER_2_1203 ();
 FILLCELL_X2 FILLER_2_1207 ();
 FILLCELL_X32 FILLER_3_1 ();
 FILLCELL_X32 FILLER_3_33 ();
 FILLCELL_X32 FILLER_3_65 ();
 FILLCELL_X32 FILLER_3_97 ();
 FILLCELL_X32 FILLER_3_129 ();
 FILLCELL_X32 FILLER_3_161 ();
 FILLCELL_X32 FILLER_3_193 ();
 FILLCELL_X32 FILLER_3_225 ();
 FILLCELL_X32 FILLER_3_257 ();
 FILLCELL_X32 FILLER_3_289 ();
 FILLCELL_X32 FILLER_3_321 ();
 FILLCELL_X32 FILLER_3_353 ();
 FILLCELL_X32 FILLER_3_385 ();
 FILLCELL_X32 FILLER_3_417 ();
 FILLCELL_X32 FILLER_3_449 ();
 FILLCELL_X32 FILLER_3_481 ();
 FILLCELL_X32 FILLER_3_513 ();
 FILLCELL_X32 FILLER_3_545 ();
 FILLCELL_X32 FILLER_3_577 ();
 FILLCELL_X4 FILLER_3_609 ();
 FILLCELL_X16 FILLER_3_650 ();
 FILLCELL_X1 FILLER_3_666 ();
 FILLCELL_X16 FILLER_3_691 ();
 FILLCELL_X1 FILLER_3_707 ();
 FILLCELL_X32 FILLER_3_734 ();
 FILLCELL_X32 FILLER_3_766 ();
 FILLCELL_X32 FILLER_3_798 ();
 FILLCELL_X32 FILLER_3_830 ();
 FILLCELL_X8 FILLER_3_862 ();
 FILLCELL_X1 FILLER_3_895 ();
 FILLCELL_X2 FILLER_3_904 ();
 FILLCELL_X2 FILLER_3_917 ();
 FILLCELL_X1 FILLER_3_919 ();
 FILLCELL_X8 FILLER_3_936 ();
 FILLCELL_X2 FILLER_3_944 ();
 FILLCELL_X4 FILLER_3_950 ();
 FILLCELL_X1 FILLER_3_954 ();
 FILLCELL_X8 FILLER_3_959 ();
 FILLCELL_X2 FILLER_3_967 ();
 FILLCELL_X8 FILLER_3_974 ();
 FILLCELL_X2 FILLER_3_982 ();
 FILLCELL_X4 FILLER_3_990 ();
 FILLCELL_X2 FILLER_3_994 ();
 FILLCELL_X1 FILLER_3_996 ();
 FILLCELL_X4 FILLER_3_1001 ();
 FILLCELL_X2 FILLER_3_1005 ();
 FILLCELL_X32 FILLER_3_1039 ();
 FILLCELL_X32 FILLER_3_1071 ();
 FILLCELL_X32 FILLER_3_1103 ();
 FILLCELL_X32 FILLER_3_1135 ();
 FILLCELL_X32 FILLER_3_1167 ();
 FILLCELL_X8 FILLER_3_1199 ();
 FILLCELL_X2 FILLER_3_1207 ();
 FILLCELL_X32 FILLER_4_1 ();
 FILLCELL_X32 FILLER_4_33 ();
 FILLCELL_X32 FILLER_4_65 ();
 FILLCELL_X32 FILLER_4_97 ();
 FILLCELL_X32 FILLER_4_129 ();
 FILLCELL_X32 FILLER_4_161 ();
 FILLCELL_X32 FILLER_4_193 ();
 FILLCELL_X32 FILLER_4_225 ();
 FILLCELL_X32 FILLER_4_257 ();
 FILLCELL_X32 FILLER_4_289 ();
 FILLCELL_X32 FILLER_4_321 ();
 FILLCELL_X8 FILLER_4_353 ();
 FILLCELL_X4 FILLER_4_361 ();
 FILLCELL_X32 FILLER_4_372 ();
 FILLCELL_X8 FILLER_4_404 ();
 FILLCELL_X2 FILLER_4_412 ();
 FILLCELL_X4 FILLER_4_423 ();
 FILLCELL_X1 FILLER_4_427 ();
 FILLCELL_X32 FILLER_4_435 ();
 FILLCELL_X32 FILLER_4_467 ();
 FILLCELL_X32 FILLER_4_499 ();
 FILLCELL_X32 FILLER_4_531 ();
 FILLCELL_X32 FILLER_4_563 ();
 FILLCELL_X16 FILLER_4_595 ();
 FILLCELL_X8 FILLER_4_611 ();
 FILLCELL_X2 FILLER_4_619 ();
 FILLCELL_X1 FILLER_4_621 ();
 FILLCELL_X2 FILLER_4_629 ();
 FILLCELL_X4 FILLER_4_632 ();
 FILLCELL_X1 FILLER_4_636 ();
 FILLCELL_X32 FILLER_4_642 ();
 FILLCELL_X32 FILLER_4_674 ();
 FILLCELL_X32 FILLER_4_706 ();
 FILLCELL_X32 FILLER_4_738 ();
 FILLCELL_X32 FILLER_4_770 ();
 FILLCELL_X32 FILLER_4_802 ();
 FILLCELL_X16 FILLER_4_834 ();
 FILLCELL_X8 FILLER_4_850 ();
 FILLCELL_X2 FILLER_4_858 ();
 FILLCELL_X8 FILLER_4_935 ();
 FILLCELL_X1 FILLER_4_943 ();
 FILLCELL_X1 FILLER_4_954 ();
 FILLCELL_X1 FILLER_4_966 ();
 FILLCELL_X4 FILLER_4_986 ();
 FILLCELL_X1 FILLER_4_990 ();
 FILLCELL_X1 FILLER_4_997 ();
 FILLCELL_X1 FILLER_4_1007 ();
 FILLCELL_X1 FILLER_4_1019 ();
 FILLCELL_X1 FILLER_4_1027 ();
 FILLCELL_X32 FILLER_4_1048 ();
 FILLCELL_X32 FILLER_4_1080 ();
 FILLCELL_X32 FILLER_4_1112 ();
 FILLCELL_X32 FILLER_4_1144 ();
 FILLCELL_X32 FILLER_4_1176 ();
 FILLCELL_X1 FILLER_4_1208 ();
 FILLCELL_X32 FILLER_5_1 ();
 FILLCELL_X32 FILLER_5_33 ();
 FILLCELL_X32 FILLER_5_65 ();
 FILLCELL_X32 FILLER_5_97 ();
 FILLCELL_X32 FILLER_5_129 ();
 FILLCELL_X32 FILLER_5_161 ();
 FILLCELL_X32 FILLER_5_193 ();
 FILLCELL_X32 FILLER_5_225 ();
 FILLCELL_X32 FILLER_5_257 ();
 FILLCELL_X32 FILLER_5_289 ();
 FILLCELL_X16 FILLER_5_321 ();
 FILLCELL_X2 FILLER_5_337 ();
 FILLCELL_X2 FILLER_5_349 ();
 FILLCELL_X1 FILLER_5_351 ();
 FILLCELL_X2 FILLER_5_362 ();
 FILLCELL_X1 FILLER_5_364 ();
 FILLCELL_X4 FILLER_5_385 ();
 FILLCELL_X2 FILLER_5_389 ();
 FILLCELL_X1 FILLER_5_391 ();
 FILLCELL_X4 FILLER_5_399 ();
 FILLCELL_X1 FILLER_5_418 ();
 FILLCELL_X1 FILLER_5_429 ();
 FILLCELL_X1 FILLER_5_437 ();
 FILLCELL_X4 FILLER_5_451 ();
 FILLCELL_X2 FILLER_5_455 ();
 FILLCELL_X1 FILLER_5_457 ();
 FILLCELL_X8 FILLER_5_483 ();
 FILLCELL_X2 FILLER_5_491 ();
 FILLCELL_X32 FILLER_5_502 ();
 FILLCELL_X32 FILLER_5_534 ();
 FILLCELL_X16 FILLER_5_566 ();
 FILLCELL_X1 FILLER_5_582 ();
 FILLCELL_X32 FILLER_5_590 ();
 FILLCELL_X32 FILLER_5_639 ();
 FILLCELL_X4 FILLER_5_671 ();
 FILLCELL_X1 FILLER_5_678 ();
 FILLCELL_X4 FILLER_5_683 ();
 FILLCELL_X1 FILLER_5_687 ();
 FILLCELL_X2 FILLER_5_692 ();
 FILLCELL_X1 FILLER_5_702 ();
 FILLCELL_X1 FILLER_5_714 ();
 FILLCELL_X32 FILLER_5_727 ();
 FILLCELL_X32 FILLER_5_759 ();
 FILLCELL_X16 FILLER_5_791 ();
 FILLCELL_X8 FILLER_5_807 ();
 FILLCELL_X2 FILLER_5_815 ();
 FILLCELL_X1 FILLER_5_817 ();
 FILLCELL_X16 FILLER_5_835 ();
 FILLCELL_X4 FILLER_5_851 ();
 FILLCELL_X2 FILLER_5_855 ();
 FILLCELL_X2 FILLER_5_874 ();
 FILLCELL_X2 FILLER_5_880 ();
 FILLCELL_X2 FILLER_5_898 ();
 FILLCELL_X8 FILLER_5_911 ();
 FILLCELL_X1 FILLER_5_919 ();
 FILLCELL_X2 FILLER_5_924 ();
 FILLCELL_X2 FILLER_5_929 ();
 FILLCELL_X8 FILLER_5_944 ();
 FILLCELL_X1 FILLER_5_952 ();
 FILLCELL_X2 FILLER_5_964 ();
 FILLCELL_X2 FILLER_5_978 ();
 FILLCELL_X1 FILLER_5_980 ();
 FILLCELL_X8 FILLER_5_986 ();
 FILLCELL_X2 FILLER_5_1012 ();
 FILLCELL_X4 FILLER_5_1037 ();
 FILLCELL_X32 FILLER_5_1048 ();
 FILLCELL_X32 FILLER_5_1080 ();
 FILLCELL_X32 FILLER_5_1112 ();
 FILLCELL_X32 FILLER_5_1144 ();
 FILLCELL_X32 FILLER_5_1176 ();
 FILLCELL_X1 FILLER_5_1208 ();
 FILLCELL_X32 FILLER_6_1 ();
 FILLCELL_X32 FILLER_6_33 ();
 FILLCELL_X32 FILLER_6_65 ();
 FILLCELL_X32 FILLER_6_97 ();
 FILLCELL_X32 FILLER_6_129 ();
 FILLCELL_X32 FILLER_6_161 ();
 FILLCELL_X32 FILLER_6_193 ();
 FILLCELL_X4 FILLER_6_225 ();
 FILLCELL_X8 FILLER_6_239 ();
 FILLCELL_X32 FILLER_6_254 ();
 FILLCELL_X32 FILLER_6_286 ();
 FILLCELL_X16 FILLER_6_318 ();
 FILLCELL_X8 FILLER_6_334 ();
 FILLCELL_X4 FILLER_6_342 ();
 FILLCELL_X2 FILLER_6_346 ();
 FILLCELL_X4 FILLER_6_353 ();
 FILLCELL_X1 FILLER_6_367 ();
 FILLCELL_X1 FILLER_6_371 ();
 FILLCELL_X1 FILLER_6_400 ();
 FILLCELL_X1 FILLER_6_412 ();
 FILLCELL_X2 FILLER_6_427 ();
 FILLCELL_X2 FILLER_6_450 ();
 FILLCELL_X1 FILLER_6_452 ();
 FILLCELL_X4 FILLER_6_460 ();
 FILLCELL_X2 FILLER_6_464 ();
 FILLCELL_X1 FILLER_6_466 ();
 FILLCELL_X32 FILLER_6_505 ();
 FILLCELL_X32 FILLER_6_537 ();
 FILLCELL_X1 FILLER_6_569 ();
 FILLCELL_X4 FILLER_6_587 ();
 FILLCELL_X4 FILLER_6_608 ();
 FILLCELL_X2 FILLER_6_612 ();
 FILLCELL_X1 FILLER_6_614 ();
 FILLCELL_X4 FILLER_6_625 ();
 FILLCELL_X2 FILLER_6_629 ();
 FILLCELL_X16 FILLER_6_632 ();
 FILLCELL_X8 FILLER_6_648 ();
 FILLCELL_X2 FILLER_6_656 ();
 FILLCELL_X2 FILLER_6_667 ();
 FILLCELL_X2 FILLER_6_690 ();
 FILLCELL_X1 FILLER_6_692 ();
 FILLCELL_X1 FILLER_6_698 ();
 FILLCELL_X1 FILLER_6_703 ();
 FILLCELL_X4 FILLER_6_708 ();
 FILLCELL_X4 FILLER_6_722 ();
 FILLCELL_X32 FILLER_6_733 ();
 FILLCELL_X32 FILLER_6_765 ();
 FILLCELL_X16 FILLER_6_797 ();
 FILLCELL_X4 FILLER_6_813 ();
 FILLCELL_X2 FILLER_6_817 ();
 FILLCELL_X1 FILLER_6_819 ();
 FILLCELL_X32 FILLER_6_827 ();
 FILLCELL_X4 FILLER_6_859 ();
 FILLCELL_X2 FILLER_6_863 ();
 FILLCELL_X1 FILLER_6_875 ();
 FILLCELL_X1 FILLER_6_888 ();
 FILLCELL_X16 FILLER_6_900 ();
 FILLCELL_X8 FILLER_6_916 ();
 FILLCELL_X4 FILLER_6_924 ();
 FILLCELL_X2 FILLER_6_928 ();
 FILLCELL_X1 FILLER_6_930 ();
 FILLCELL_X1 FILLER_6_941 ();
 FILLCELL_X4 FILLER_6_946 ();
 FILLCELL_X2 FILLER_6_950 ();
 FILLCELL_X4 FILLER_6_959 ();
 FILLCELL_X2 FILLER_6_975 ();
 FILLCELL_X4 FILLER_6_981 ();
 FILLCELL_X1 FILLER_6_990 ();
 FILLCELL_X2 FILLER_6_1040 ();
 FILLCELL_X1 FILLER_6_1042 ();
 FILLCELL_X32 FILLER_6_1050 ();
 FILLCELL_X32 FILLER_6_1082 ();
 FILLCELL_X32 FILLER_6_1114 ();
 FILLCELL_X32 FILLER_6_1146 ();
 FILLCELL_X16 FILLER_6_1178 ();
 FILLCELL_X8 FILLER_6_1194 ();
 FILLCELL_X4 FILLER_6_1202 ();
 FILLCELL_X2 FILLER_6_1206 ();
 FILLCELL_X1 FILLER_6_1208 ();
 FILLCELL_X32 FILLER_7_1 ();
 FILLCELL_X32 FILLER_7_33 ();
 FILLCELL_X32 FILLER_7_65 ();
 FILLCELL_X32 FILLER_7_97 ();
 FILLCELL_X32 FILLER_7_129 ();
 FILLCELL_X16 FILLER_7_161 ();
 FILLCELL_X8 FILLER_7_190 ();
 FILLCELL_X4 FILLER_7_198 ();
 FILLCELL_X8 FILLER_7_209 ();
 FILLCELL_X1 FILLER_7_217 ();
 FILLCELL_X4 FILLER_7_230 ();
 FILLCELL_X2 FILLER_7_234 ();
 FILLCELL_X1 FILLER_7_236 ();
 FILLCELL_X2 FILLER_7_250 ();
 FILLCELL_X1 FILLER_7_252 ();
 FILLCELL_X32 FILLER_7_289 ();
 FILLCELL_X16 FILLER_7_321 ();
 FILLCELL_X8 FILLER_7_337 ();
 FILLCELL_X1 FILLER_7_345 ();
 FILLCELL_X4 FILLER_7_356 ();
 FILLCELL_X2 FILLER_7_360 ();
 FILLCELL_X1 FILLER_7_362 ();
 FILLCELL_X1 FILLER_7_375 ();
 FILLCELL_X2 FILLER_7_400 ();
 FILLCELL_X1 FILLER_7_402 ();
 FILLCELL_X2 FILLER_7_418 ();
 FILLCELL_X2 FILLER_7_469 ();
 FILLCELL_X1 FILLER_7_471 ();
 FILLCELL_X32 FILLER_7_498 ();
 FILLCELL_X32 FILLER_7_530 ();
 FILLCELL_X32 FILLER_7_562 ();
 FILLCELL_X4 FILLER_7_594 ();
 FILLCELL_X1 FILLER_7_611 ();
 FILLCELL_X8 FILLER_7_643 ();
 FILLCELL_X4 FILLER_7_651 ();
 FILLCELL_X2 FILLER_7_659 ();
 FILLCELL_X1 FILLER_7_661 ();
 FILLCELL_X1 FILLER_7_665 ();
 FILLCELL_X8 FILLER_7_671 ();
 FILLCELL_X4 FILLER_7_679 ();
 FILLCELL_X1 FILLER_7_683 ();
 FILLCELL_X4 FILLER_7_690 ();
 FILLCELL_X1 FILLER_7_694 ();
 FILLCELL_X1 FILLER_7_705 ();
 FILLCELL_X2 FILLER_7_717 ();
 FILLCELL_X8 FILLER_7_726 ();
 FILLCELL_X4 FILLER_7_741 ();
 FILLCELL_X2 FILLER_7_745 ();
 FILLCELL_X32 FILLER_7_759 ();
 FILLCELL_X16 FILLER_7_791 ();
 FILLCELL_X8 FILLER_7_807 ();
 FILLCELL_X4 FILLER_7_815 ();
 FILLCELL_X2 FILLER_7_819 ();
 FILLCELL_X1 FILLER_7_821 ();
 FILLCELL_X16 FILLER_7_839 ();
 FILLCELL_X8 FILLER_7_855 ();
 FILLCELL_X4 FILLER_7_863 ();
 FILLCELL_X4 FILLER_7_871 ();
 FILLCELL_X8 FILLER_7_878 ();
 FILLCELL_X1 FILLER_7_886 ();
 FILLCELL_X4 FILLER_7_905 ();
 FILLCELL_X1 FILLER_7_913 ();
 FILLCELL_X4 FILLER_7_920 ();
 FILLCELL_X1 FILLER_7_924 ();
 FILLCELL_X8 FILLER_7_928 ();
 FILLCELL_X4 FILLER_7_936 ();
 FILLCELL_X2 FILLER_7_940 ();
 FILLCELL_X2 FILLER_7_949 ();
 FILLCELL_X4 FILLER_7_960 ();
 FILLCELL_X2 FILLER_7_964 ();
 FILLCELL_X8 FILLER_7_977 ();
 FILLCELL_X4 FILLER_7_985 ();
 FILLCELL_X2 FILLER_7_989 ();
 FILLCELL_X1 FILLER_7_991 ();
 FILLCELL_X8 FILLER_7_999 ();
 FILLCELL_X2 FILLER_7_1007 ();
 FILLCELL_X2 FILLER_7_1029 ();
 FILLCELL_X4 FILLER_7_1041 ();
 FILLCELL_X1 FILLER_7_1045 ();
 FILLCELL_X32 FILLER_7_1068 ();
 FILLCELL_X32 FILLER_7_1100 ();
 FILLCELL_X32 FILLER_7_1132 ();
 FILLCELL_X32 FILLER_7_1164 ();
 FILLCELL_X8 FILLER_7_1196 ();
 FILLCELL_X4 FILLER_7_1204 ();
 FILLCELL_X1 FILLER_7_1208 ();
 FILLCELL_X32 FILLER_8_1 ();
 FILLCELL_X32 FILLER_8_33 ();
 FILLCELL_X32 FILLER_8_65 ();
 FILLCELL_X32 FILLER_8_97 ();
 FILLCELL_X32 FILLER_8_129 ();
 FILLCELL_X2 FILLER_8_161 ();
 FILLCELL_X1 FILLER_8_163 ();
 FILLCELL_X1 FILLER_8_223 ();
 FILLCELL_X1 FILLER_8_233 ();
 FILLCELL_X1 FILLER_8_241 ();
 FILLCELL_X2 FILLER_8_255 ();
 FILLCELL_X32 FILLER_8_302 ();
 FILLCELL_X8 FILLER_8_334 ();
 FILLCELL_X4 FILLER_8_342 ();
 FILLCELL_X2 FILLER_8_346 ();
 FILLCELL_X1 FILLER_8_348 ();
 FILLCELL_X4 FILLER_8_362 ();
 FILLCELL_X2 FILLER_8_386 ();
 FILLCELL_X1 FILLER_8_388 ();
 FILLCELL_X1 FILLER_8_396 ();
 FILLCELL_X1 FILLER_8_404 ();
 FILLCELL_X1 FILLER_8_412 ();
 FILLCELL_X1 FILLER_8_420 ();
 FILLCELL_X4 FILLER_8_445 ();
 FILLCELL_X2 FILLER_8_449 ();
 FILLCELL_X1 FILLER_8_451 ();
 FILLCELL_X2 FILLER_8_454 ();
 FILLCELL_X1 FILLER_8_456 ();
 FILLCELL_X2 FILLER_8_464 ();
 FILLCELL_X2 FILLER_8_473 ();
 FILLCELL_X2 FILLER_8_482 ();
 FILLCELL_X1 FILLER_8_484 ();
 FILLCELL_X32 FILLER_8_493 ();
 FILLCELL_X32 FILLER_8_525 ();
 FILLCELL_X16 FILLER_8_557 ();
 FILLCELL_X8 FILLER_8_573 ();
 FILLCELL_X4 FILLER_8_581 ();
 FILLCELL_X8 FILLER_8_602 ();
 FILLCELL_X2 FILLER_8_610 ();
 FILLCELL_X1 FILLER_8_612 ();
 FILLCELL_X8 FILLER_8_616 ();
 FILLCELL_X2 FILLER_8_629 ();
 FILLCELL_X16 FILLER_8_632 ();
 FILLCELL_X8 FILLER_8_648 ();
 FILLCELL_X4 FILLER_8_656 ();
 FILLCELL_X2 FILLER_8_660 ();
 FILLCELL_X1 FILLER_8_662 ();
 FILLCELL_X1 FILLER_8_667 ();
 FILLCELL_X4 FILLER_8_685 ();
 FILLCELL_X1 FILLER_8_689 ();
 FILLCELL_X16 FILLER_8_697 ();
 FILLCELL_X2 FILLER_8_713 ();
 FILLCELL_X1 FILLER_8_715 ();
 FILLCELL_X4 FILLER_8_719 ();
 FILLCELL_X2 FILLER_8_739 ();
 FILLCELL_X1 FILLER_8_741 ();
 FILLCELL_X32 FILLER_8_756 ();
 FILLCELL_X32 FILLER_8_788 ();
 FILLCELL_X16 FILLER_8_820 ();
 FILLCELL_X8 FILLER_8_836 ();
 FILLCELL_X4 FILLER_8_844 ();
 FILLCELL_X2 FILLER_8_848 ();
 FILLCELL_X4 FILLER_8_867 ();
 FILLCELL_X2 FILLER_8_871 ();
 FILLCELL_X1 FILLER_8_873 ();
 FILLCELL_X2 FILLER_8_900 ();
 FILLCELL_X2 FILLER_8_913 ();
 FILLCELL_X1 FILLER_8_915 ();
 FILLCELL_X1 FILLER_8_920 ();
 FILLCELL_X4 FILLER_8_925 ();
 FILLCELL_X2 FILLER_8_937 ();
 FILLCELL_X1 FILLER_8_939 ();
 FILLCELL_X4 FILLER_8_948 ();
 FILLCELL_X4 FILLER_8_970 ();
 FILLCELL_X1 FILLER_8_974 ();
 FILLCELL_X2 FILLER_8_989 ();
 FILLCELL_X2 FILLER_8_997 ();
 FILLCELL_X1 FILLER_8_999 ();
 FILLCELL_X2 FILLER_8_1005 ();
 FILLCELL_X16 FILLER_8_1022 ();
 FILLCELL_X1 FILLER_8_1057 ();
 FILLCELL_X32 FILLER_8_1065 ();
 FILLCELL_X32 FILLER_8_1097 ();
 FILLCELL_X32 FILLER_8_1129 ();
 FILLCELL_X32 FILLER_8_1161 ();
 FILLCELL_X16 FILLER_8_1193 ();
 FILLCELL_X32 FILLER_9_1 ();
 FILLCELL_X32 FILLER_9_33 ();
 FILLCELL_X32 FILLER_9_65 ();
 FILLCELL_X32 FILLER_9_97 ();
 FILLCELL_X32 FILLER_9_129 ();
 FILLCELL_X4 FILLER_9_161 ();
 FILLCELL_X2 FILLER_9_165 ();
 FILLCELL_X2 FILLER_9_171 ();
 FILLCELL_X4 FILLER_9_179 ();
 FILLCELL_X2 FILLER_9_183 ();
 FILLCELL_X2 FILLER_9_240 ();
 FILLCELL_X2 FILLER_9_265 ();
 FILLCELL_X2 FILLER_9_274 ();
 FILLCELL_X1 FILLER_9_276 ();
 FILLCELL_X32 FILLER_9_296 ();
 FILLCELL_X16 FILLER_9_328 ();
 FILLCELL_X4 FILLER_9_344 ();
 FILLCELL_X1 FILLER_9_362 ();
 FILLCELL_X4 FILLER_9_403 ();
 FILLCELL_X1 FILLER_9_417 ();
 FILLCELL_X4 FILLER_9_447 ();
 FILLCELL_X2 FILLER_9_468 ();
 FILLCELL_X32 FILLER_9_489 ();
 FILLCELL_X32 FILLER_9_521 ();
 FILLCELL_X32 FILLER_9_553 ();
 FILLCELL_X16 FILLER_9_585 ();
 FILLCELL_X4 FILLER_9_601 ();
 FILLCELL_X4 FILLER_9_612 ();
 FILLCELL_X2 FILLER_9_641 ();
 FILLCELL_X2 FILLER_9_654 ();
 FILLCELL_X2 FILLER_9_670 ();
 FILLCELL_X1 FILLER_9_672 ();
 FILLCELL_X2 FILLER_9_688 ();
 FILLCELL_X1 FILLER_9_690 ();
 FILLCELL_X4 FILLER_9_697 ();
 FILLCELL_X4 FILLER_9_712 ();
 FILLCELL_X2 FILLER_9_716 ();
 FILLCELL_X2 FILLER_9_735 ();
 FILLCELL_X1 FILLER_9_737 ();
 FILLCELL_X32 FILLER_9_763 ();
 FILLCELL_X16 FILLER_9_795 ();
 FILLCELL_X8 FILLER_9_811 ();
 FILLCELL_X32 FILLER_9_824 ();
 FILLCELL_X8 FILLER_9_856 ();
 FILLCELL_X2 FILLER_9_864 ();
 FILLCELL_X1 FILLER_9_866 ();
 FILLCELL_X4 FILLER_9_873 ();
 FILLCELL_X1 FILLER_9_877 ();
 FILLCELL_X4 FILLER_9_886 ();
 FILLCELL_X1 FILLER_9_890 ();
 FILLCELL_X2 FILLER_9_905 ();
 FILLCELL_X1 FILLER_9_907 ();
 FILLCELL_X4 FILLER_9_911 ();
 FILLCELL_X16 FILLER_9_931 ();
 FILLCELL_X1 FILLER_9_947 ();
 FILLCELL_X2 FILLER_9_951 ();
 FILLCELL_X1 FILLER_9_953 ();
 FILLCELL_X1 FILLER_9_957 ();
 FILLCELL_X1 FILLER_9_962 ();
 FILLCELL_X1 FILLER_9_986 ();
 FILLCELL_X4 FILLER_9_1002 ();
 FILLCELL_X4 FILLER_9_1009 ();
 FILLCELL_X2 FILLER_9_1017 ();
 FILLCELL_X2 FILLER_9_1030 ();
 FILLCELL_X1 FILLER_9_1032 ();
 FILLCELL_X4 FILLER_9_1044 ();
 FILLCELL_X2 FILLER_9_1048 ();
 FILLCELL_X1 FILLER_9_1050 ();
 FILLCELL_X1 FILLER_9_1054 ();
 FILLCELL_X32 FILLER_9_1065 ();
 FILLCELL_X32 FILLER_9_1097 ();
 FILLCELL_X32 FILLER_9_1129 ();
 FILLCELL_X32 FILLER_9_1161 ();
 FILLCELL_X16 FILLER_9_1193 ();
 FILLCELL_X32 FILLER_10_1 ();
 FILLCELL_X32 FILLER_10_33 ();
 FILLCELL_X32 FILLER_10_65 ();
 FILLCELL_X32 FILLER_10_97 ();
 FILLCELL_X32 FILLER_10_129 ();
 FILLCELL_X2 FILLER_10_161 ();
 FILLCELL_X1 FILLER_10_171 ();
 FILLCELL_X4 FILLER_10_182 ();
 FILLCELL_X1 FILLER_10_186 ();
 FILLCELL_X8 FILLER_10_194 ();
 FILLCELL_X1 FILLER_10_220 ();
 FILLCELL_X4 FILLER_10_267 ();
 FILLCELL_X2 FILLER_10_271 ();
 FILLCELL_X4 FILLER_10_280 ();
 FILLCELL_X32 FILLER_10_307 ();
 FILLCELL_X16 FILLER_10_339 ();
 FILLCELL_X1 FILLER_10_355 ();
 FILLCELL_X2 FILLER_10_366 ();
 FILLCELL_X2 FILLER_10_414 ();
 FILLCELL_X16 FILLER_10_423 ();
 FILLCELL_X2 FILLER_10_446 ();
 FILLCELL_X4 FILLER_10_458 ();
 FILLCELL_X32 FILLER_10_502 ();
 FILLCELL_X32 FILLER_10_534 ();
 FILLCELL_X2 FILLER_10_566 ();
 FILLCELL_X1 FILLER_10_578 ();
 FILLCELL_X2 FILLER_10_584 ();
 FILLCELL_X1 FILLER_10_586 ();
 FILLCELL_X4 FILLER_10_613 ();
 FILLCELL_X2 FILLER_10_617 ();
 FILLCELL_X1 FILLER_10_619 ();
 FILLCELL_X1 FILLER_10_624 ();
 FILLCELL_X2 FILLER_10_629 ();
 FILLCELL_X1 FILLER_10_648 ();
 FILLCELL_X1 FILLER_10_662 ();
 FILLCELL_X2 FILLER_10_671 ();
 FILLCELL_X2 FILLER_10_682 ();
 FILLCELL_X4 FILLER_10_695 ();
 FILLCELL_X2 FILLER_10_699 ();
 FILLCELL_X4 FILLER_10_720 ();
 FILLCELL_X4 FILLER_10_729 ();
 FILLCELL_X2 FILLER_10_733 ();
 FILLCELL_X2 FILLER_10_748 ();
 FILLCELL_X32 FILLER_10_761 ();
 FILLCELL_X32 FILLER_10_793 ();
 FILLCELL_X8 FILLER_10_825 ();
 FILLCELL_X1 FILLER_10_833 ();
 FILLCELL_X16 FILLER_10_841 ();
 FILLCELL_X8 FILLER_10_857 ();
 FILLCELL_X4 FILLER_10_865 ();
 FILLCELL_X2 FILLER_10_869 ();
 FILLCELL_X1 FILLER_10_877 ();
 FILLCELL_X4 FILLER_10_897 ();
 FILLCELL_X1 FILLER_10_901 ();
 FILLCELL_X1 FILLER_10_910 ();
 FILLCELL_X1 FILLER_10_918 ();
 FILLCELL_X1 FILLER_10_925 ();
 FILLCELL_X1 FILLER_10_936 ();
 FILLCELL_X4 FILLER_10_948 ();
 FILLCELL_X2 FILLER_10_952 ();
 FILLCELL_X8 FILLER_10_957 ();
 FILLCELL_X2 FILLER_10_965 ();
 FILLCELL_X1 FILLER_10_967 ();
 FILLCELL_X4 FILLER_10_975 ();
 FILLCELL_X1 FILLER_10_979 ();
 FILLCELL_X4 FILLER_10_1009 ();
 FILLCELL_X1 FILLER_10_1013 ();
 FILLCELL_X2 FILLER_10_1017 ();
 FILLCELL_X1 FILLER_10_1019 ();
 FILLCELL_X2 FILLER_10_1023 ();
 FILLCELL_X1 FILLER_10_1041 ();
 FILLCELL_X32 FILLER_10_1057 ();
 FILLCELL_X32 FILLER_10_1089 ();
 FILLCELL_X32 FILLER_10_1121 ();
 FILLCELL_X32 FILLER_10_1153 ();
 FILLCELL_X16 FILLER_10_1185 ();
 FILLCELL_X8 FILLER_10_1201 ();
 FILLCELL_X32 FILLER_11_1 ();
 FILLCELL_X32 FILLER_11_33 ();
 FILLCELL_X32 FILLER_11_65 ();
 FILLCELL_X32 FILLER_11_97 ();
 FILLCELL_X4 FILLER_11_129 ();
 FILLCELL_X2 FILLER_11_133 ();
 FILLCELL_X1 FILLER_11_135 ();
 FILLCELL_X8 FILLER_11_146 ();
 FILLCELL_X1 FILLER_11_165 ();
 FILLCELL_X2 FILLER_11_188 ();
 FILLCELL_X4 FILLER_11_210 ();
 FILLCELL_X1 FILLER_11_221 ();
 FILLCELL_X4 FILLER_11_277 ();
 FILLCELL_X2 FILLER_11_281 ();
 FILLCELL_X1 FILLER_11_296 ();
 FILLCELL_X32 FILLER_11_311 ();
 FILLCELL_X2 FILLER_11_343 ();
 FILLCELL_X1 FILLER_11_358 ();
 FILLCELL_X1 FILLER_11_384 ();
 FILLCELL_X2 FILLER_11_392 ();
 FILLCELL_X2 FILLER_11_401 ();
 FILLCELL_X16 FILLER_11_425 ();
 FILLCELL_X1 FILLER_11_441 ();
 FILLCELL_X4 FILLER_11_463 ();
 FILLCELL_X2 FILLER_11_467 ();
 FILLCELL_X2 FILLER_11_488 ();
 FILLCELL_X1 FILLER_11_490 ();
 FILLCELL_X32 FILLER_11_500 ();
 FILLCELL_X32 FILLER_11_532 ();
 FILLCELL_X16 FILLER_11_564 ();
 FILLCELL_X8 FILLER_11_598 ();
 FILLCELL_X1 FILLER_11_606 ();
 FILLCELL_X8 FILLER_11_614 ();
 FILLCELL_X2 FILLER_11_627 ();
 FILLCELL_X8 FILLER_11_633 ();
 FILLCELL_X1 FILLER_11_641 ();
 FILLCELL_X1 FILLER_11_667 ();
 FILLCELL_X4 FILLER_11_701 ();
 FILLCELL_X2 FILLER_11_705 ();
 FILLCELL_X1 FILLER_11_707 ();
 FILLCELL_X4 FILLER_11_716 ();
 FILLCELL_X4 FILLER_11_728 ();
 FILLCELL_X1 FILLER_11_732 ();
 FILLCELL_X1 FILLER_11_737 ();
 FILLCELL_X4 FILLER_11_760 ();
 FILLCELL_X32 FILLER_11_775 ();
 FILLCELL_X32 FILLER_11_807 ();
 FILLCELL_X16 FILLER_11_839 ();
 FILLCELL_X8 FILLER_11_855 ();
 FILLCELL_X4 FILLER_11_863 ();
 FILLCELL_X2 FILLER_11_867 ();
 FILLCELL_X1 FILLER_11_869 ();
 FILLCELL_X1 FILLER_11_886 ();
 FILLCELL_X1 FILLER_11_896 ();
 FILLCELL_X4 FILLER_11_900 ();
 FILLCELL_X2 FILLER_11_904 ();
 FILLCELL_X1 FILLER_11_906 ();
 FILLCELL_X2 FILLER_11_912 ();
 FILLCELL_X1 FILLER_11_914 ();
 FILLCELL_X2 FILLER_11_922 ();
 FILLCELL_X2 FILLER_11_935 ();
 FILLCELL_X1 FILLER_11_937 ();
 FILLCELL_X1 FILLER_11_941 ();
 FILLCELL_X4 FILLER_11_953 ();
 FILLCELL_X1 FILLER_11_957 ();
 FILLCELL_X2 FILLER_11_983 ();
 FILLCELL_X1 FILLER_11_997 ();
 FILLCELL_X2 FILLER_11_1012 ();
 FILLCELL_X1 FILLER_11_1014 ();
 FILLCELL_X2 FILLER_11_1019 ();
 FILLCELL_X2 FILLER_11_1035 ();
 FILLCELL_X32 FILLER_11_1054 ();
 FILLCELL_X32 FILLER_11_1086 ();
 FILLCELL_X32 FILLER_11_1118 ();
 FILLCELL_X32 FILLER_11_1150 ();
 FILLCELL_X16 FILLER_11_1182 ();
 FILLCELL_X8 FILLER_11_1198 ();
 FILLCELL_X2 FILLER_11_1206 ();
 FILLCELL_X1 FILLER_11_1208 ();
 FILLCELL_X32 FILLER_12_1 ();
 FILLCELL_X32 FILLER_12_33 ();
 FILLCELL_X32 FILLER_12_65 ();
 FILLCELL_X32 FILLER_12_97 ();
 FILLCELL_X8 FILLER_12_129 ();
 FILLCELL_X4 FILLER_12_137 ();
 FILLCELL_X2 FILLER_12_146 ();
 FILLCELL_X1 FILLER_12_148 ();
 FILLCELL_X4 FILLER_12_153 ();
 FILLCELL_X2 FILLER_12_157 ();
 FILLCELL_X2 FILLER_12_171 ();
 FILLCELL_X1 FILLER_12_173 ();
 FILLCELL_X1 FILLER_12_192 ();
 FILLCELL_X2 FILLER_12_196 ();
 FILLCELL_X1 FILLER_12_198 ();
 FILLCELL_X4 FILLER_12_211 ();
 FILLCELL_X1 FILLER_12_228 ();
 FILLCELL_X4 FILLER_12_235 ();
 FILLCELL_X32 FILLER_12_313 ();
 FILLCELL_X8 FILLER_12_345 ();
 FILLCELL_X1 FILLER_12_353 ();
 FILLCELL_X1 FILLER_12_376 ();
 FILLCELL_X2 FILLER_12_394 ();
 FILLCELL_X2 FILLER_12_425 ();
 FILLCELL_X1 FILLER_12_427 ();
 FILLCELL_X2 FILLER_12_430 ();
 FILLCELL_X2 FILLER_12_441 ();
 FILLCELL_X1 FILLER_12_443 ();
 FILLCELL_X1 FILLER_12_451 ();
 FILLCELL_X4 FILLER_12_459 ();
 FILLCELL_X1 FILLER_12_463 ();
 FILLCELL_X2 FILLER_12_474 ();
 FILLCELL_X1 FILLER_12_483 ();
 FILLCELL_X2 FILLER_12_491 ();
 FILLCELL_X1 FILLER_12_493 ();
 FILLCELL_X32 FILLER_12_501 ();
 FILLCELL_X32 FILLER_12_533 ();
 FILLCELL_X32 FILLER_12_565 ();
 FILLCELL_X1 FILLER_12_597 ();
 FILLCELL_X1 FILLER_12_616 ();
 FILLCELL_X4 FILLER_12_650 ();
 FILLCELL_X2 FILLER_12_654 ();
 FILLCELL_X1 FILLER_12_686 ();
 FILLCELL_X1 FILLER_12_702 ();
 FILLCELL_X2 FILLER_12_715 ();
 FILLCELL_X1 FILLER_12_717 ();
 FILLCELL_X4 FILLER_12_722 ();
 FILLCELL_X2 FILLER_12_726 ();
 FILLCELL_X1 FILLER_12_728 ();
 FILLCELL_X1 FILLER_12_747 ();
 FILLCELL_X1 FILLER_12_758 ();
 FILLCELL_X32 FILLER_12_767 ();
 FILLCELL_X32 FILLER_12_799 ();
 FILLCELL_X32 FILLER_12_831 ();
 FILLCELL_X4 FILLER_12_863 ();
 FILLCELL_X2 FILLER_12_867 ();
 FILLCELL_X1 FILLER_12_869 ();
 FILLCELL_X2 FILLER_12_873 ();
 FILLCELL_X1 FILLER_12_875 ();
 FILLCELL_X2 FILLER_12_893 ();
 FILLCELL_X1 FILLER_12_895 ();
 FILLCELL_X2 FILLER_12_899 ();
 FILLCELL_X4 FILLER_12_910 ();
 FILLCELL_X1 FILLER_12_914 ();
 FILLCELL_X1 FILLER_12_918 ();
 FILLCELL_X1 FILLER_12_926 ();
 FILLCELL_X8 FILLER_12_940 ();
 FILLCELL_X2 FILLER_12_948 ();
 FILLCELL_X1 FILLER_12_950 ();
 FILLCELL_X2 FILLER_12_956 ();
 FILLCELL_X2 FILLER_12_962 ();
 FILLCELL_X4 FILLER_12_968 ();
 FILLCELL_X2 FILLER_12_972 ();
 FILLCELL_X1 FILLER_12_974 ();
 FILLCELL_X1 FILLER_12_982 ();
 FILLCELL_X2 FILLER_12_1005 ();
 FILLCELL_X1 FILLER_12_1034 ();
 FILLCELL_X32 FILLER_12_1042 ();
 FILLCELL_X32 FILLER_12_1074 ();
 FILLCELL_X32 FILLER_12_1106 ();
 FILLCELL_X32 FILLER_12_1138 ();
 FILLCELL_X32 FILLER_12_1170 ();
 FILLCELL_X4 FILLER_12_1202 ();
 FILLCELL_X2 FILLER_12_1206 ();
 FILLCELL_X1 FILLER_12_1208 ();
 FILLCELL_X32 FILLER_13_1 ();
 FILLCELL_X32 FILLER_13_33 ();
 FILLCELL_X32 FILLER_13_65 ();
 FILLCELL_X32 FILLER_13_97 ();
 FILLCELL_X8 FILLER_13_129 ();
 FILLCELL_X2 FILLER_13_137 ();
 FILLCELL_X1 FILLER_13_139 ();
 FILLCELL_X4 FILLER_13_150 ();
 FILLCELL_X2 FILLER_13_154 ();
 FILLCELL_X1 FILLER_13_156 ();
 FILLCELL_X2 FILLER_13_178 ();
 FILLCELL_X1 FILLER_13_180 ();
 FILLCELL_X2 FILLER_13_186 ();
 FILLCELL_X1 FILLER_13_191 ();
 FILLCELL_X8 FILLER_13_200 ();
 FILLCELL_X2 FILLER_13_208 ();
 FILLCELL_X1 FILLER_13_214 ();
 FILLCELL_X2 FILLER_13_222 ();
 FILLCELL_X2 FILLER_13_239 ();
 FILLCELL_X2 FILLER_13_253 ();
 FILLCELL_X2 FILLER_13_288 ();
 FILLCELL_X4 FILLER_13_297 ();
 FILLCELL_X16 FILLER_13_308 ();
 FILLCELL_X8 FILLER_13_324 ();
 FILLCELL_X2 FILLER_13_332 ();
 FILLCELL_X1 FILLER_13_334 ();
 FILLCELL_X8 FILLER_13_344 ();
 FILLCELL_X2 FILLER_13_352 ();
 FILLCELL_X1 FILLER_13_354 ();
 FILLCELL_X2 FILLER_13_370 ();
 FILLCELL_X1 FILLER_13_414 ();
 FILLCELL_X1 FILLER_13_419 ();
 FILLCELL_X4 FILLER_13_430 ();
 FILLCELL_X2 FILLER_13_434 ();
 FILLCELL_X4 FILLER_13_445 ();
 FILLCELL_X2 FILLER_13_449 ();
 FILLCELL_X1 FILLER_13_451 ();
 FILLCELL_X2 FILLER_13_491 ();
 FILLCELL_X32 FILLER_13_505 ();
 FILLCELL_X32 FILLER_13_537 ();
 FILLCELL_X8 FILLER_13_569 ();
 FILLCELL_X2 FILLER_13_615 ();
 FILLCELL_X4 FILLER_13_626 ();
 FILLCELL_X8 FILLER_13_655 ();
 FILLCELL_X16 FILLER_13_704 ();
 FILLCELL_X8 FILLER_13_720 ();
 FILLCELL_X4 FILLER_13_728 ();
 FILLCELL_X8 FILLER_13_736 ();
 FILLCELL_X2 FILLER_13_747 ();
 FILLCELL_X1 FILLER_13_749 ();
 FILLCELL_X2 FILLER_13_754 ();
 FILLCELL_X1 FILLER_13_756 ();
 FILLCELL_X4 FILLER_13_769 ();
 FILLCELL_X32 FILLER_13_798 ();
 FILLCELL_X16 FILLER_13_830 ();
 FILLCELL_X4 FILLER_13_846 ();
 FILLCELL_X1 FILLER_13_850 ();
 FILLCELL_X4 FILLER_13_863 ();
 FILLCELL_X1 FILLER_13_885 ();
 FILLCELL_X8 FILLER_13_908 ();
 FILLCELL_X2 FILLER_13_916 ();
 FILLCELL_X4 FILLER_13_925 ();
 FILLCELL_X2 FILLER_13_929 ();
 FILLCELL_X8 FILLER_13_937 ();
 FILLCELL_X4 FILLER_13_945 ();
 FILLCELL_X2 FILLER_13_949 ();
 FILLCELL_X8 FILLER_13_963 ();
 FILLCELL_X2 FILLER_13_971 ();
 FILLCELL_X1 FILLER_13_973 ();
 FILLCELL_X4 FILLER_13_986 ();
 FILLCELL_X2 FILLER_13_1002 ();
 FILLCELL_X1 FILLER_13_1004 ();
 FILLCELL_X2 FILLER_13_1012 ();
 FILLCELL_X1 FILLER_13_1014 ();
 FILLCELL_X4 FILLER_13_1018 ();
 FILLCELL_X2 FILLER_13_1022 ();
 FILLCELL_X32 FILLER_13_1048 ();
 FILLCELL_X32 FILLER_13_1080 ();
 FILLCELL_X32 FILLER_13_1112 ();
 FILLCELL_X32 FILLER_13_1144 ();
 FILLCELL_X32 FILLER_13_1176 ();
 FILLCELL_X1 FILLER_13_1208 ();
 FILLCELL_X32 FILLER_14_1 ();
 FILLCELL_X32 FILLER_14_33 ();
 FILLCELL_X32 FILLER_14_65 ();
 FILLCELL_X32 FILLER_14_97 ();
 FILLCELL_X16 FILLER_14_129 ();
 FILLCELL_X4 FILLER_14_145 ();
 FILLCELL_X2 FILLER_14_149 ();
 FILLCELL_X2 FILLER_14_170 ();
 FILLCELL_X2 FILLER_14_183 ();
 FILLCELL_X2 FILLER_14_192 ();
 FILLCELL_X1 FILLER_14_198 ();
 FILLCELL_X4 FILLER_14_202 ();
 FILLCELL_X1 FILLER_14_222 ();
 FILLCELL_X1 FILLER_14_231 ();
 FILLCELL_X4 FILLER_14_237 ();
 FILLCELL_X1 FILLER_14_241 ();
 FILLCELL_X2 FILLER_14_257 ();
 FILLCELL_X4 FILLER_14_304 ();
 FILLCELL_X2 FILLER_14_308 ();
 FILLCELL_X16 FILLER_14_319 ();
 FILLCELL_X4 FILLER_14_335 ();
 FILLCELL_X1 FILLER_14_339 ();
 FILLCELL_X1 FILLER_14_385 ();
 FILLCELL_X1 FILLER_14_407 ();
 FILLCELL_X1 FILLER_14_432 ();
 FILLCELL_X8 FILLER_14_447 ();
 FILLCELL_X2 FILLER_14_455 ();
 FILLCELL_X1 FILLER_14_457 ();
 FILLCELL_X4 FILLER_14_462 ();
 FILLCELL_X1 FILLER_14_466 ();
 FILLCELL_X2 FILLER_14_480 ();
 FILLCELL_X1 FILLER_14_482 ();
 FILLCELL_X32 FILLER_14_501 ();
 FILLCELL_X32 FILLER_14_533 ();
 FILLCELL_X32 FILLER_14_565 ();
 FILLCELL_X2 FILLER_14_597 ();
 FILLCELL_X1 FILLER_14_599 ();
 FILLCELL_X1 FILLER_14_615 ();
 FILLCELL_X1 FILLER_14_625 ();
 FILLCELL_X1 FILLER_14_639 ();
 FILLCELL_X1 FILLER_14_647 ();
 FILLCELL_X1 FILLER_14_664 ();
 FILLCELL_X8 FILLER_14_679 ();
 FILLCELL_X1 FILLER_14_687 ();
 FILLCELL_X2 FILLER_14_692 ();
 FILLCELL_X1 FILLER_14_694 ();
 FILLCELL_X4 FILLER_14_710 ();
 FILLCELL_X1 FILLER_14_720 ();
 FILLCELL_X4 FILLER_14_729 ();
 FILLCELL_X1 FILLER_14_733 ();
 FILLCELL_X1 FILLER_14_739 ();
 FILLCELL_X2 FILLER_14_743 ();
 FILLCELL_X32 FILLER_14_766 ();
 FILLCELL_X32 FILLER_14_798 ();
 FILLCELL_X32 FILLER_14_830 ();
 FILLCELL_X4 FILLER_14_862 ();
 FILLCELL_X2 FILLER_14_866 ();
 FILLCELL_X1 FILLER_14_875 ();
 FILLCELL_X2 FILLER_14_894 ();
 FILLCELL_X1 FILLER_14_896 ();
 FILLCELL_X8 FILLER_14_903 ();
 FILLCELL_X4 FILLER_14_911 ();
 FILLCELL_X2 FILLER_14_915 ();
 FILLCELL_X1 FILLER_14_917 ();
 FILLCELL_X1 FILLER_14_925 ();
 FILLCELL_X4 FILLER_14_944 ();
 FILLCELL_X2 FILLER_14_948 ();
 FILLCELL_X1 FILLER_14_962 ();
 FILLCELL_X2 FILLER_14_973 ();
 FILLCELL_X4 FILLER_14_1008 ();
 FILLCELL_X32 FILLER_14_1055 ();
 FILLCELL_X32 FILLER_14_1087 ();
 FILLCELL_X32 FILLER_14_1119 ();
 FILLCELL_X32 FILLER_14_1151 ();
 FILLCELL_X16 FILLER_14_1183 ();
 FILLCELL_X8 FILLER_14_1199 ();
 FILLCELL_X2 FILLER_14_1207 ();
 FILLCELL_X32 FILLER_15_1 ();
 FILLCELL_X32 FILLER_15_33 ();
 FILLCELL_X32 FILLER_15_65 ();
 FILLCELL_X32 FILLER_15_97 ();
 FILLCELL_X32 FILLER_15_129 ();
 FILLCELL_X16 FILLER_15_161 ();
 FILLCELL_X2 FILLER_15_177 ();
 FILLCELL_X4 FILLER_15_194 ();
 FILLCELL_X16 FILLER_15_210 ();
 FILLCELL_X2 FILLER_15_226 ();
 FILLCELL_X1 FILLER_15_247 ();
 FILLCELL_X1 FILLER_15_255 ();
 FILLCELL_X2 FILLER_15_263 ();
 FILLCELL_X1 FILLER_15_265 ();
 FILLCELL_X1 FILLER_15_293 ();
 FILLCELL_X32 FILLER_15_307 ();
 FILLCELL_X8 FILLER_15_339 ();
 FILLCELL_X4 FILLER_15_347 ();
 FILLCELL_X2 FILLER_15_377 ();
 FILLCELL_X4 FILLER_15_386 ();
 FILLCELL_X2 FILLER_15_390 ();
 FILLCELL_X8 FILLER_15_400 ();
 FILLCELL_X4 FILLER_15_408 ();
 FILLCELL_X2 FILLER_15_420 ();
 FILLCELL_X1 FILLER_15_422 ();
 FILLCELL_X4 FILLER_15_454 ();
 FILLCELL_X2 FILLER_15_458 ();
 FILLCELL_X2 FILLER_15_474 ();
 FILLCELL_X16 FILLER_15_499 ();
 FILLCELL_X8 FILLER_15_515 ();
 FILLCELL_X4 FILLER_15_523 ();
 FILLCELL_X2 FILLER_15_527 ();
 FILLCELL_X1 FILLER_15_529 ();
 FILLCELL_X16 FILLER_15_537 ();
 FILLCELL_X8 FILLER_15_553 ();
 FILLCELL_X1 FILLER_15_561 ();
 FILLCELL_X16 FILLER_15_579 ();
 FILLCELL_X2 FILLER_15_595 ();
 FILLCELL_X1 FILLER_15_597 ();
 FILLCELL_X2 FILLER_15_609 ();
 FILLCELL_X2 FILLER_15_615 ();
 FILLCELL_X1 FILLER_15_617 ();
 FILLCELL_X2 FILLER_15_623 ();
 FILLCELL_X8 FILLER_15_629 ();
 FILLCELL_X1 FILLER_15_668 ();
 FILLCELL_X2 FILLER_15_680 ();
 FILLCELL_X2 FILLER_15_684 ();
 FILLCELL_X4 FILLER_15_690 ();
 FILLCELL_X1 FILLER_15_694 ();
 FILLCELL_X4 FILLER_15_715 ();
 FILLCELL_X2 FILLER_15_719 ();
 FILLCELL_X1 FILLER_15_721 ();
 FILLCELL_X32 FILLER_15_759 ();
 FILLCELL_X32 FILLER_15_791 ();
 FILLCELL_X32 FILLER_15_823 ();
 FILLCELL_X16 FILLER_15_855 ();
 FILLCELL_X1 FILLER_15_871 ();
 FILLCELL_X1 FILLER_15_875 ();
 FILLCELL_X2 FILLER_15_880 ();
 FILLCELL_X1 FILLER_15_882 ();
 FILLCELL_X8 FILLER_15_897 ();
 FILLCELL_X1 FILLER_15_926 ();
 FILLCELL_X4 FILLER_15_932 ();
 FILLCELL_X8 FILLER_15_940 ();
 FILLCELL_X4 FILLER_15_948 ();
 FILLCELL_X2 FILLER_15_952 ();
 FILLCELL_X1 FILLER_15_963 ();
 FILLCELL_X1 FILLER_15_971 ();
 FILLCELL_X4 FILLER_15_976 ();
 FILLCELL_X2 FILLER_15_987 ();
 FILLCELL_X1 FILLER_15_989 ();
 FILLCELL_X2 FILLER_15_1001 ();
 FILLCELL_X1 FILLER_15_1003 ();
 FILLCELL_X1 FILLER_15_1010 ();
 FILLCELL_X2 FILLER_15_1016 ();
 FILLCELL_X2 FILLER_15_1032 ();
 FILLCELL_X32 FILLER_15_1056 ();
 FILLCELL_X32 FILLER_15_1088 ();
 FILLCELL_X32 FILLER_15_1120 ();
 FILLCELL_X32 FILLER_15_1152 ();
 FILLCELL_X16 FILLER_15_1184 ();
 FILLCELL_X8 FILLER_15_1200 ();
 FILLCELL_X1 FILLER_15_1208 ();
 FILLCELL_X32 FILLER_16_1 ();
 FILLCELL_X32 FILLER_16_33 ();
 FILLCELL_X32 FILLER_16_65 ();
 FILLCELL_X32 FILLER_16_97 ();
 FILLCELL_X8 FILLER_16_129 ();
 FILLCELL_X4 FILLER_16_137 ();
 FILLCELL_X2 FILLER_16_141 ();
 FILLCELL_X1 FILLER_16_143 ();
 FILLCELL_X2 FILLER_16_153 ();
 FILLCELL_X1 FILLER_16_155 ();
 FILLCELL_X1 FILLER_16_186 ();
 FILLCELL_X4 FILLER_16_198 ();
 FILLCELL_X2 FILLER_16_202 ();
 FILLCELL_X2 FILLER_16_208 ();
 FILLCELL_X1 FILLER_16_210 ();
 FILLCELL_X1 FILLER_16_219 ();
 FILLCELL_X1 FILLER_16_223 ();
 FILLCELL_X4 FILLER_16_232 ();
 FILLCELL_X1 FILLER_16_236 ();
 FILLCELL_X1 FILLER_16_280 ();
 FILLCELL_X32 FILLER_16_306 ();
 FILLCELL_X8 FILLER_16_338 ();
 FILLCELL_X1 FILLER_16_346 ();
 FILLCELL_X1 FILLER_16_365 ();
 FILLCELL_X2 FILLER_16_373 ();
 FILLCELL_X1 FILLER_16_379 ();
 FILLCELL_X2 FILLER_16_386 ();
 FILLCELL_X1 FILLER_16_393 ();
 FILLCELL_X1 FILLER_16_425 ();
 FILLCELL_X2 FILLER_16_429 ();
 FILLCELL_X2 FILLER_16_442 ();
 FILLCELL_X4 FILLER_16_457 ();
 FILLCELL_X2 FILLER_16_461 ();
 FILLCELL_X4 FILLER_16_486 ();
 FILLCELL_X1 FILLER_16_490 ();
 FILLCELL_X16 FILLER_16_498 ();
 FILLCELL_X4 FILLER_16_514 ();
 FILLCELL_X1 FILLER_16_518 ();
 FILLCELL_X32 FILLER_16_538 ();
 FILLCELL_X4 FILLER_16_570 ();
 FILLCELL_X2 FILLER_16_574 ();
 FILLCELL_X1 FILLER_16_576 ();
 FILLCELL_X4 FILLER_16_587 ();
 FILLCELL_X1 FILLER_16_591 ();
 FILLCELL_X2 FILLER_16_607 ();
 FILLCELL_X1 FILLER_16_609 ();
 FILLCELL_X2 FILLER_16_628 ();
 FILLCELL_X1 FILLER_16_630 ();
 FILLCELL_X2 FILLER_16_649 ();
 FILLCELL_X1 FILLER_16_651 ();
 FILLCELL_X2 FILLER_16_687 ();
 FILLCELL_X4 FILLER_16_694 ();
 FILLCELL_X2 FILLER_16_703 ();
 FILLCELL_X1 FILLER_16_705 ();
 FILLCELL_X2 FILLER_16_718 ();
 FILLCELL_X1 FILLER_16_720 ();
 FILLCELL_X2 FILLER_16_724 ();
 FILLCELL_X1 FILLER_16_726 ();
 FILLCELL_X16 FILLER_16_731 ();
 FILLCELL_X2 FILLER_16_747 ();
 FILLCELL_X8 FILLER_16_761 ();
 FILLCELL_X1 FILLER_16_769 ();
 FILLCELL_X8 FILLER_16_787 ();
 FILLCELL_X32 FILLER_16_812 ();
 FILLCELL_X16 FILLER_16_844 ();
 FILLCELL_X1 FILLER_16_860 ();
 FILLCELL_X2 FILLER_16_868 ();
 FILLCELL_X1 FILLER_16_870 ();
 FILLCELL_X1 FILLER_16_889 ();
 FILLCELL_X2 FILLER_16_909 ();
 FILLCELL_X2 FILLER_16_925 ();
 FILLCELL_X4 FILLER_16_938 ();
 FILLCELL_X1 FILLER_16_942 ();
 FILLCELL_X8 FILLER_16_948 ();
 FILLCELL_X1 FILLER_16_956 ();
 FILLCELL_X8 FILLER_16_961 ();
 FILLCELL_X2 FILLER_16_979 ();
 FILLCELL_X1 FILLER_16_1002 ();
 FILLCELL_X2 FILLER_16_1009 ();
 FILLCELL_X2 FILLER_16_1014 ();
 FILLCELL_X1 FILLER_16_1016 ();
 FILLCELL_X4 FILLER_16_1031 ();
 FILLCELL_X2 FILLER_16_1035 ();
 FILLCELL_X1 FILLER_16_1037 ();
 FILLCELL_X1 FILLER_16_1052 ();
 FILLCELL_X32 FILLER_16_1056 ();
 FILLCELL_X32 FILLER_16_1088 ();
 FILLCELL_X32 FILLER_16_1120 ();
 FILLCELL_X32 FILLER_16_1152 ();
 FILLCELL_X16 FILLER_16_1184 ();
 FILLCELL_X8 FILLER_16_1200 ();
 FILLCELL_X1 FILLER_16_1208 ();
 FILLCELL_X32 FILLER_17_1 ();
 FILLCELL_X32 FILLER_17_33 ();
 FILLCELL_X32 FILLER_17_65 ();
 FILLCELL_X32 FILLER_17_97 ();
 FILLCELL_X4 FILLER_17_129 ();
 FILLCELL_X2 FILLER_17_133 ();
 FILLCELL_X4 FILLER_17_139 ();
 FILLCELL_X2 FILLER_17_148 ();
 FILLCELL_X1 FILLER_17_150 ();
 FILLCELL_X4 FILLER_17_154 ();
 FILLCELL_X1 FILLER_17_158 ();
 FILLCELL_X2 FILLER_17_177 ();
 FILLCELL_X1 FILLER_17_179 ();
 FILLCELL_X4 FILLER_17_191 ();
 FILLCELL_X1 FILLER_17_195 ();
 FILLCELL_X2 FILLER_17_212 ();
 FILLCELL_X4 FILLER_17_225 ();
 FILLCELL_X2 FILLER_17_235 ();
 FILLCELL_X1 FILLER_17_278 ();
 FILLCELL_X2 FILLER_17_292 ();
 FILLCELL_X32 FILLER_17_297 ();
 FILLCELL_X8 FILLER_17_329 ();
 FILLCELL_X4 FILLER_17_337 ();
 FILLCELL_X1 FILLER_17_341 ();
 FILLCELL_X1 FILLER_17_353 ();
 FILLCELL_X8 FILLER_17_365 ();
 FILLCELL_X4 FILLER_17_373 ();
 FILLCELL_X1 FILLER_17_384 ();
 FILLCELL_X1 FILLER_17_389 ();
 FILLCELL_X1 FILLER_17_397 ();
 FILLCELL_X1 FILLER_17_403 ();
 FILLCELL_X2 FILLER_17_415 ();
 FILLCELL_X1 FILLER_17_417 ();
 FILLCELL_X4 FILLER_17_421 ();
 FILLCELL_X1 FILLER_17_428 ();
 FILLCELL_X4 FILLER_17_434 ();
 FILLCELL_X1 FILLER_17_444 ();
 FILLCELL_X2 FILLER_17_467 ();
 FILLCELL_X32 FILLER_17_500 ();
 FILLCELL_X32 FILLER_17_532 ();
 FILLCELL_X4 FILLER_17_564 ();
 FILLCELL_X2 FILLER_17_568 ();
 FILLCELL_X4 FILLER_17_587 ();
 FILLCELL_X2 FILLER_17_591 ();
 FILLCELL_X1 FILLER_17_593 ();
 FILLCELL_X8 FILLER_17_597 ();
 FILLCELL_X1 FILLER_17_605 ();
 FILLCELL_X1 FILLER_17_609 ();
 FILLCELL_X1 FILLER_17_613 ();
 FILLCELL_X4 FILLER_17_632 ();
 FILLCELL_X1 FILLER_17_636 ();
 FILLCELL_X4 FILLER_17_652 ();
 FILLCELL_X2 FILLER_17_656 ();
 FILLCELL_X2 FILLER_17_669 ();
 FILLCELL_X1 FILLER_17_676 ();
 FILLCELL_X8 FILLER_17_687 ();
 FILLCELL_X1 FILLER_17_695 ();
 FILLCELL_X2 FILLER_17_707 ();
 FILLCELL_X4 FILLER_17_714 ();
 FILLCELL_X2 FILLER_17_718 ();
 FILLCELL_X8 FILLER_17_723 ();
 FILLCELL_X2 FILLER_17_731 ();
 FILLCELL_X1 FILLER_17_733 ();
 FILLCELL_X2 FILLER_17_746 ();
 FILLCELL_X1 FILLER_17_748 ();
 FILLCELL_X1 FILLER_17_753 ();
 FILLCELL_X16 FILLER_17_757 ();
 FILLCELL_X2 FILLER_17_773 ();
 FILLCELL_X1 FILLER_17_775 ();
 FILLCELL_X32 FILLER_17_783 ();
 FILLCELL_X32 FILLER_17_815 ();
 FILLCELL_X8 FILLER_17_847 ();
 FILLCELL_X2 FILLER_17_855 ();
 FILLCELL_X1 FILLER_17_857 ();
 FILLCELL_X2 FILLER_17_879 ();
 FILLCELL_X2 FILLER_17_885 ();
 FILLCELL_X2 FILLER_17_911 ();
 FILLCELL_X1 FILLER_17_913 ();
 FILLCELL_X2 FILLER_17_930 ();
 FILLCELL_X1 FILLER_17_932 ();
 FILLCELL_X4 FILLER_17_952 ();
 FILLCELL_X2 FILLER_17_956 ();
 FILLCELL_X1 FILLER_17_958 ();
 FILLCELL_X1 FILLER_17_967 ();
 FILLCELL_X1 FILLER_17_971 ();
 FILLCELL_X2 FILLER_17_992 ();
 FILLCELL_X1 FILLER_17_994 ();
 FILLCELL_X4 FILLER_17_1021 ();
 FILLCELL_X2 FILLER_17_1047 ();
 FILLCELL_X32 FILLER_17_1053 ();
 FILLCELL_X32 FILLER_17_1085 ();
 FILLCELL_X32 FILLER_17_1117 ();
 FILLCELL_X32 FILLER_17_1149 ();
 FILLCELL_X16 FILLER_17_1181 ();
 FILLCELL_X8 FILLER_17_1197 ();
 FILLCELL_X4 FILLER_17_1205 ();
 FILLCELL_X32 FILLER_18_1 ();
 FILLCELL_X32 FILLER_18_33 ();
 FILLCELL_X32 FILLER_18_65 ();
 FILLCELL_X32 FILLER_18_97 ();
 FILLCELL_X1 FILLER_18_129 ();
 FILLCELL_X4 FILLER_18_134 ();
 FILLCELL_X2 FILLER_18_138 ();
 FILLCELL_X2 FILLER_18_155 ();
 FILLCELL_X1 FILLER_18_157 ();
 FILLCELL_X2 FILLER_18_196 ();
 FILLCELL_X4 FILLER_18_214 ();
 FILLCELL_X8 FILLER_18_229 ();
 FILLCELL_X4 FILLER_18_237 ();
 FILLCELL_X1 FILLER_18_258 ();
 FILLCELL_X2 FILLER_18_297 ();
 FILLCELL_X1 FILLER_18_299 ();
 FILLCELL_X16 FILLER_18_313 ();
 FILLCELL_X2 FILLER_18_329 ();
 FILLCELL_X1 FILLER_18_331 ();
 FILLCELL_X2 FILLER_18_352 ();
 FILLCELL_X1 FILLER_18_357 ();
 FILLCELL_X1 FILLER_18_365 ();
 FILLCELL_X2 FILLER_18_378 ();
 FILLCELL_X1 FILLER_18_380 ();
 FILLCELL_X1 FILLER_18_388 ();
 FILLCELL_X2 FILLER_18_396 ();
 FILLCELL_X1 FILLER_18_398 ();
 FILLCELL_X4 FILLER_18_402 ();
 FILLCELL_X2 FILLER_18_406 ();
 FILLCELL_X2 FILLER_18_412 ();
 FILLCELL_X1 FILLER_18_418 ();
 FILLCELL_X4 FILLER_18_427 ();
 FILLCELL_X2 FILLER_18_431 ();
 FILLCELL_X1 FILLER_18_433 ();
 FILLCELL_X4 FILLER_18_446 ();
 FILLCELL_X2 FILLER_18_454 ();
 FILLCELL_X8 FILLER_18_461 ();
 FILLCELL_X1 FILLER_18_469 ();
 FILLCELL_X1 FILLER_18_488 ();
 FILLCELL_X32 FILLER_18_500 ();
 FILLCELL_X32 FILLER_18_532 ();
 FILLCELL_X2 FILLER_18_564 ();
 FILLCELL_X1 FILLER_18_566 ();
 FILLCELL_X4 FILLER_18_584 ();
 FILLCELL_X1 FILLER_18_588 ();
 FILLCELL_X2 FILLER_18_602 ();
 FILLCELL_X1 FILLER_18_604 ();
 FILLCELL_X2 FILLER_18_620 ();
 FILLCELL_X1 FILLER_18_622 ();
 FILLCELL_X4 FILLER_18_632 ();
 FILLCELL_X2 FILLER_18_636 ();
 FILLCELL_X1 FILLER_18_638 ();
 FILLCELL_X8 FILLER_18_646 ();
 FILLCELL_X8 FILLER_18_690 ();
 FILLCELL_X2 FILLER_18_698 ();
 FILLCELL_X1 FILLER_18_700 ();
 FILLCELL_X1 FILLER_18_707 ();
 FILLCELL_X2 FILLER_18_715 ();
 FILLCELL_X1 FILLER_18_721 ();
 FILLCELL_X4 FILLER_18_726 ();
 FILLCELL_X2 FILLER_18_734 ();
 FILLCELL_X1 FILLER_18_736 ();
 FILLCELL_X32 FILLER_18_751 ();
 FILLCELL_X32 FILLER_18_783 ();
 FILLCELL_X32 FILLER_18_815 ();
 FILLCELL_X8 FILLER_18_847 ();
 FILLCELL_X1 FILLER_18_874 ();
 FILLCELL_X2 FILLER_18_881 ();
 FILLCELL_X2 FILLER_18_898 ();
 FILLCELL_X1 FILLER_18_900 ();
 FILLCELL_X1 FILLER_18_904 ();
 FILLCELL_X2 FILLER_18_927 ();
 FILLCELL_X4 FILLER_18_940 ();
 FILLCELL_X4 FILLER_18_949 ();
 FILLCELL_X1 FILLER_18_953 ();
 FILLCELL_X1 FILLER_18_987 ();
 FILLCELL_X1 FILLER_18_1001 ();
 FILLCELL_X2 FILLER_18_1019 ();
 FILLCELL_X1 FILLER_18_1028 ();
 FILLCELL_X32 FILLER_18_1049 ();
 FILLCELL_X32 FILLER_18_1081 ();
 FILLCELL_X32 FILLER_18_1113 ();
 FILLCELL_X32 FILLER_18_1145 ();
 FILLCELL_X32 FILLER_18_1177 ();
 FILLCELL_X32 FILLER_19_1 ();
 FILLCELL_X32 FILLER_19_33 ();
 FILLCELL_X32 FILLER_19_65 ();
 FILLCELL_X16 FILLER_19_97 ();
 FILLCELL_X8 FILLER_19_113 ();
 FILLCELL_X4 FILLER_19_121 ();
 FILLCELL_X2 FILLER_19_125 ();
 FILLCELL_X1 FILLER_19_138 ();
 FILLCELL_X1 FILLER_19_155 ();
 FILLCELL_X1 FILLER_19_190 ();
 FILLCELL_X4 FILLER_19_201 ();
 FILLCELL_X1 FILLER_19_205 ();
 FILLCELL_X1 FILLER_19_222 ();
 FILLCELL_X32 FILLER_19_305 ();
 FILLCELL_X8 FILLER_19_337 ();
 FILLCELL_X4 FILLER_19_379 ();
 FILLCELL_X2 FILLER_19_383 ();
 FILLCELL_X1 FILLER_19_403 ();
 FILLCELL_X8 FILLER_19_412 ();
 FILLCELL_X2 FILLER_19_420 ();
 FILLCELL_X1 FILLER_19_446 ();
 FILLCELL_X1 FILLER_19_450 ();
 FILLCELL_X2 FILLER_19_463 ();
 FILLCELL_X1 FILLER_19_465 ();
 FILLCELL_X32 FILLER_19_494 ();
 FILLCELL_X16 FILLER_19_526 ();
 FILLCELL_X2 FILLER_19_542 ();
 FILLCELL_X1 FILLER_19_544 ();
 FILLCELL_X4 FILLER_19_560 ();
 FILLCELL_X1 FILLER_19_564 ();
 FILLCELL_X8 FILLER_19_589 ();
 FILLCELL_X1 FILLER_19_597 ();
 FILLCELL_X2 FILLER_19_607 ();
 FILLCELL_X1 FILLER_19_609 ();
 FILLCELL_X16 FILLER_19_618 ();
 FILLCELL_X4 FILLER_19_634 ();
 FILLCELL_X2 FILLER_19_652 ();
 FILLCELL_X1 FILLER_19_654 ();
 FILLCELL_X8 FILLER_19_662 ();
 FILLCELL_X4 FILLER_19_670 ();
 FILLCELL_X1 FILLER_19_674 ();
 FILLCELL_X4 FILLER_19_680 ();
 FILLCELL_X2 FILLER_19_684 ();
 FILLCELL_X1 FILLER_19_686 ();
 FILLCELL_X8 FILLER_19_698 ();
 FILLCELL_X2 FILLER_19_706 ();
 FILLCELL_X1 FILLER_19_708 ();
 FILLCELL_X4 FILLER_19_714 ();
 FILLCELL_X1 FILLER_19_718 ();
 FILLCELL_X1 FILLER_19_728 ();
 FILLCELL_X2 FILLER_19_747 ();
 FILLCELL_X1 FILLER_19_749 ();
 FILLCELL_X1 FILLER_19_763 ();
 FILLCELL_X32 FILLER_19_774 ();
 FILLCELL_X8 FILLER_19_806 ();
 FILLCELL_X16 FILLER_19_821 ();
 FILLCELL_X4 FILLER_19_837 ();
 FILLCELL_X2 FILLER_19_841 ();
 FILLCELL_X2 FILLER_19_860 ();
 FILLCELL_X1 FILLER_19_862 ();
 FILLCELL_X1 FILLER_19_874 ();
 FILLCELL_X4 FILLER_19_878 ();
 FILLCELL_X1 FILLER_19_882 ();
 FILLCELL_X2 FILLER_19_902 ();
 FILLCELL_X2 FILLER_19_908 ();
 FILLCELL_X1 FILLER_19_910 ();
 FILLCELL_X4 FILLER_19_922 ();
 FILLCELL_X2 FILLER_19_933 ();
 FILLCELL_X2 FILLER_19_946 ();
 FILLCELL_X1 FILLER_19_977 ();
 FILLCELL_X1 FILLER_19_987 ();
 FILLCELL_X2 FILLER_19_1029 ();
 FILLCELL_X8 FILLER_19_1041 ();
 FILLCELL_X2 FILLER_19_1049 ();
 FILLCELL_X32 FILLER_19_1065 ();
 FILLCELL_X32 FILLER_19_1097 ();
 FILLCELL_X32 FILLER_19_1129 ();
 FILLCELL_X32 FILLER_19_1161 ();
 FILLCELL_X16 FILLER_19_1193 ();
 FILLCELL_X32 FILLER_20_1 ();
 FILLCELL_X32 FILLER_20_33 ();
 FILLCELL_X32 FILLER_20_65 ();
 FILLCELL_X16 FILLER_20_97 ();
 FILLCELL_X8 FILLER_20_113 ();
 FILLCELL_X4 FILLER_20_121 ();
 FILLCELL_X1 FILLER_20_125 ();
 FILLCELL_X1 FILLER_20_135 ();
 FILLCELL_X16 FILLER_20_160 ();
 FILLCELL_X8 FILLER_20_176 ();
 FILLCELL_X4 FILLER_20_184 ();
 FILLCELL_X1 FILLER_20_214 ();
 FILLCELL_X4 FILLER_20_222 ();
 FILLCELL_X2 FILLER_20_244 ();
 FILLCELL_X2 FILLER_20_251 ();
 FILLCELL_X2 FILLER_20_275 ();
 FILLCELL_X1 FILLER_20_292 ();
 FILLCELL_X16 FILLER_20_312 ();
 FILLCELL_X4 FILLER_20_328 ();
 FILLCELL_X4 FILLER_20_339 ();
 FILLCELL_X2 FILLER_20_343 ();
 FILLCELL_X1 FILLER_20_354 ();
 FILLCELL_X1 FILLER_20_361 ();
 FILLCELL_X2 FILLER_20_365 ();
 FILLCELL_X4 FILLER_20_374 ();
 FILLCELL_X2 FILLER_20_378 ();
 FILLCELL_X1 FILLER_20_384 ();
 FILLCELL_X16 FILLER_20_392 ();
 FILLCELL_X2 FILLER_20_408 ();
 FILLCELL_X1 FILLER_20_410 ();
 FILLCELL_X4 FILLER_20_427 ();
 FILLCELL_X2 FILLER_20_431 ();
 FILLCELL_X4 FILLER_20_437 ();
 FILLCELL_X2 FILLER_20_444 ();
 FILLCELL_X4 FILLER_20_494 ();
 FILLCELL_X2 FILLER_20_498 ();
 FILLCELL_X16 FILLER_20_503 ();
 FILLCELL_X4 FILLER_20_519 ();
 FILLCELL_X2 FILLER_20_523 ();
 FILLCELL_X1 FILLER_20_525 ();
 FILLCELL_X2 FILLER_20_562 ();
 FILLCELL_X4 FILLER_20_613 ();
 FILLCELL_X2 FILLER_20_617 ();
 FILLCELL_X2 FILLER_20_632 ();
 FILLCELL_X1 FILLER_20_634 ();
 FILLCELL_X4 FILLER_20_646 ();
 FILLCELL_X2 FILLER_20_671 ();
 FILLCELL_X1 FILLER_20_673 ();
 FILLCELL_X4 FILLER_20_678 ();
 FILLCELL_X1 FILLER_20_682 ();
 FILLCELL_X4 FILLER_20_686 ();
 FILLCELL_X2 FILLER_20_690 ();
 FILLCELL_X1 FILLER_20_692 ();
 FILLCELL_X2 FILLER_20_701 ();
 FILLCELL_X1 FILLER_20_703 ();
 FILLCELL_X4 FILLER_20_708 ();
 FILLCELL_X4 FILLER_20_714 ();
 FILLCELL_X2 FILLER_20_718 ();
 FILLCELL_X1 FILLER_20_720 ();
 FILLCELL_X2 FILLER_20_725 ();
 FILLCELL_X2 FILLER_20_731 ();
 FILLCELL_X2 FILLER_20_752 ();
 FILLCELL_X2 FILLER_20_761 ();
 FILLCELL_X32 FILLER_20_765 ();
 FILLCELL_X32 FILLER_20_797 ();
 FILLCELL_X32 FILLER_20_829 ();
 FILLCELL_X16 FILLER_20_861 ();
 FILLCELL_X2 FILLER_20_877 ();
 FILLCELL_X1 FILLER_20_879 ();
 FILLCELL_X1 FILLER_20_895 ();
 FILLCELL_X4 FILLER_20_907 ();
 FILLCELL_X2 FILLER_20_916 ();
 FILLCELL_X2 FILLER_20_922 ();
 FILLCELL_X1 FILLER_20_926 ();
 FILLCELL_X2 FILLER_20_934 ();
 FILLCELL_X1 FILLER_20_957 ();
 FILLCELL_X2 FILLER_20_991 ();
 FILLCELL_X2 FILLER_20_1034 ();
 FILLCELL_X1 FILLER_20_1036 ();
 FILLCELL_X32 FILLER_20_1060 ();
 FILLCELL_X32 FILLER_20_1092 ();
 FILLCELL_X32 FILLER_20_1124 ();
 FILLCELL_X32 FILLER_20_1156 ();
 FILLCELL_X16 FILLER_20_1188 ();
 FILLCELL_X4 FILLER_20_1204 ();
 FILLCELL_X1 FILLER_20_1208 ();
 FILLCELL_X32 FILLER_21_1 ();
 FILLCELL_X32 FILLER_21_33 ();
 FILLCELL_X32 FILLER_21_65 ();
 FILLCELL_X16 FILLER_21_97 ();
 FILLCELL_X8 FILLER_21_113 ();
 FILLCELL_X4 FILLER_21_121 ();
 FILLCELL_X2 FILLER_21_125 ();
 FILLCELL_X2 FILLER_21_134 ();
 FILLCELL_X1 FILLER_21_136 ();
 FILLCELL_X1 FILLER_21_144 ();
 FILLCELL_X1 FILLER_21_156 ();
 FILLCELL_X2 FILLER_21_168 ();
 FILLCELL_X2 FILLER_21_173 ();
 FILLCELL_X4 FILLER_21_181 ();
 FILLCELL_X2 FILLER_21_185 ();
 FILLCELL_X1 FILLER_21_187 ();
 FILLCELL_X8 FILLER_21_199 ();
 FILLCELL_X2 FILLER_21_207 ();
 FILLCELL_X1 FILLER_21_209 ();
 FILLCELL_X1 FILLER_21_216 ();
 FILLCELL_X2 FILLER_21_278 ();
 FILLCELL_X1 FILLER_21_280 ();
 FILLCELL_X2 FILLER_21_286 ();
 FILLCELL_X1 FILLER_21_288 ();
 FILLCELL_X1 FILLER_21_301 ();
 FILLCELL_X2 FILLER_21_316 ();
 FILLCELL_X4 FILLER_21_337 ();
 FILLCELL_X2 FILLER_21_355 ();
 FILLCELL_X1 FILLER_21_360 ();
 FILLCELL_X1 FILLER_21_372 ();
 FILLCELL_X1 FILLER_21_380 ();
 FILLCELL_X2 FILLER_21_385 ();
 FILLCELL_X1 FILLER_21_387 ();
 FILLCELL_X1 FILLER_21_393 ();
 FILLCELL_X4 FILLER_21_396 ();
 FILLCELL_X2 FILLER_21_400 ();
 FILLCELL_X2 FILLER_21_409 ();
 FILLCELL_X1 FILLER_21_411 ();
 FILLCELL_X2 FILLER_21_416 ();
 FILLCELL_X1 FILLER_21_418 ();
 FILLCELL_X4 FILLER_21_428 ();
 FILLCELL_X1 FILLER_21_432 ();
 FILLCELL_X2 FILLER_21_437 ();
 FILLCELL_X1 FILLER_21_439 ();
 FILLCELL_X2 FILLER_21_445 ();
 FILLCELL_X4 FILLER_21_451 ();
 FILLCELL_X2 FILLER_21_463 ();
 FILLCELL_X32 FILLER_21_490 ();
 FILLCELL_X16 FILLER_21_522 ();
 FILLCELL_X4 FILLER_21_538 ();
 FILLCELL_X2 FILLER_21_549 ();
 FILLCELL_X1 FILLER_21_551 ();
 FILLCELL_X8 FILLER_21_578 ();
 FILLCELL_X4 FILLER_21_612 ();
 FILLCELL_X2 FILLER_21_616 ();
 FILLCELL_X1 FILLER_21_618 ();
 FILLCELL_X2 FILLER_21_626 ();
 FILLCELL_X1 FILLER_21_632 ();
 FILLCELL_X2 FILLER_21_642 ();
 FILLCELL_X1 FILLER_21_659 ();
 FILLCELL_X4 FILLER_21_665 ();
 FILLCELL_X1 FILLER_21_669 ();
 FILLCELL_X4 FILLER_21_673 ();
 FILLCELL_X2 FILLER_21_696 ();
 FILLCELL_X2 FILLER_21_705 ();
 FILLCELL_X2 FILLER_21_736 ();
 FILLCELL_X1 FILLER_21_738 ();
 FILLCELL_X32 FILLER_21_742 ();
 FILLCELL_X16 FILLER_21_774 ();
 FILLCELL_X8 FILLER_21_790 ();
 FILLCELL_X1 FILLER_21_798 ();
 FILLCELL_X32 FILLER_21_816 ();
 FILLCELL_X32 FILLER_21_848 ();
 FILLCELL_X4 FILLER_21_880 ();
 FILLCELL_X2 FILLER_21_884 ();
 FILLCELL_X1 FILLER_21_886 ();
 FILLCELL_X2 FILLER_21_900 ();
 FILLCELL_X1 FILLER_21_902 ();
 FILLCELL_X4 FILLER_21_912 ();
 FILLCELL_X1 FILLER_21_916 ();
 FILLCELL_X1 FILLER_21_954 ();
 FILLCELL_X2 FILLER_21_1022 ();
 FILLCELL_X32 FILLER_21_1055 ();
 FILLCELL_X32 FILLER_21_1087 ();
 FILLCELL_X32 FILLER_21_1119 ();
 FILLCELL_X32 FILLER_21_1151 ();
 FILLCELL_X16 FILLER_21_1183 ();
 FILLCELL_X8 FILLER_21_1199 ();
 FILLCELL_X2 FILLER_21_1207 ();
 FILLCELL_X32 FILLER_22_1 ();
 FILLCELL_X32 FILLER_22_33 ();
 FILLCELL_X32 FILLER_22_65 ();
 FILLCELL_X16 FILLER_22_97 ();
 FILLCELL_X8 FILLER_22_113 ();
 FILLCELL_X2 FILLER_22_121 ();
 FILLCELL_X1 FILLER_22_123 ();
 FILLCELL_X2 FILLER_22_142 ();
 FILLCELL_X1 FILLER_22_144 ();
 FILLCELL_X4 FILLER_22_156 ();
 FILLCELL_X2 FILLER_22_227 ();
 FILLCELL_X1 FILLER_22_265 ();
 FILLCELL_X2 FILLER_22_273 ();
 FILLCELL_X32 FILLER_22_305 ();
 FILLCELL_X2 FILLER_22_337 ();
 FILLCELL_X4 FILLER_22_344 ();
 FILLCELL_X2 FILLER_22_355 ();
 FILLCELL_X1 FILLER_22_357 ();
 FILLCELL_X8 FILLER_22_368 ();
 FILLCELL_X2 FILLER_22_376 ();
 FILLCELL_X2 FILLER_22_389 ();
 FILLCELL_X1 FILLER_22_391 ();
 FILLCELL_X2 FILLER_22_402 ();
 FILLCELL_X2 FILLER_22_408 ();
 FILLCELL_X1 FILLER_22_410 ();
 FILLCELL_X4 FILLER_22_418 ();
 FILLCELL_X1 FILLER_22_422 ();
 FILLCELL_X4 FILLER_22_454 ();
 FILLCELL_X1 FILLER_22_458 ();
 FILLCELL_X2 FILLER_22_464 ();
 FILLCELL_X1 FILLER_22_466 ();
 FILLCELL_X32 FILLER_22_491 ();
 FILLCELL_X8 FILLER_22_523 ();
 FILLCELL_X1 FILLER_22_531 ();
 FILLCELL_X8 FILLER_22_568 ();
 FILLCELL_X4 FILLER_22_576 ();
 FILLCELL_X2 FILLER_22_596 ();
 FILLCELL_X1 FILLER_22_598 ();
 FILLCELL_X4 FILLER_22_612 ();
 FILLCELL_X1 FILLER_22_616 ();
 FILLCELL_X2 FILLER_22_622 ();
 FILLCELL_X1 FILLER_22_639 ();
 FILLCELL_X2 FILLER_22_649 ();
 FILLCELL_X1 FILLER_22_651 ();
 FILLCELL_X16 FILLER_22_660 ();
 FILLCELL_X2 FILLER_22_676 ();
 FILLCELL_X1 FILLER_22_678 ();
 FILLCELL_X4 FILLER_22_687 ();
 FILLCELL_X2 FILLER_22_691 ();
 FILLCELL_X16 FILLER_22_702 ();
 FILLCELL_X8 FILLER_22_718 ();
 FILLCELL_X1 FILLER_22_726 ();
 FILLCELL_X8 FILLER_22_741 ();
 FILLCELL_X2 FILLER_22_749 ();
 FILLCELL_X16 FILLER_22_762 ();
 FILLCELL_X8 FILLER_22_778 ();
 FILLCELL_X2 FILLER_22_786 ();
 FILLCELL_X1 FILLER_22_834 ();
 FILLCELL_X8 FILLER_22_854 ();
 FILLCELL_X1 FILLER_22_878 ();
 FILLCELL_X8 FILLER_22_886 ();
 FILLCELL_X2 FILLER_22_894 ();
 FILLCELL_X1 FILLER_22_896 ();
 FILLCELL_X4 FILLER_22_906 ();
 FILLCELL_X4 FILLER_22_923 ();
 FILLCELL_X1 FILLER_22_927 ();
 FILLCELL_X8 FILLER_22_942 ();
 FILLCELL_X2 FILLER_22_969 ();
 FILLCELL_X1 FILLER_22_982 ();
 FILLCELL_X32 FILLER_22_1041 ();
 FILLCELL_X32 FILLER_22_1073 ();
 FILLCELL_X32 FILLER_22_1105 ();
 FILLCELL_X32 FILLER_22_1137 ();
 FILLCELL_X32 FILLER_22_1169 ();
 FILLCELL_X8 FILLER_22_1201 ();
 FILLCELL_X32 FILLER_23_1 ();
 FILLCELL_X32 FILLER_23_33 ();
 FILLCELL_X32 FILLER_23_65 ();
 FILLCELL_X16 FILLER_23_97 ();
 FILLCELL_X8 FILLER_23_113 ();
 FILLCELL_X2 FILLER_23_121 ();
 FILLCELL_X2 FILLER_23_134 ();
 FILLCELL_X1 FILLER_23_136 ();
 FILLCELL_X2 FILLER_23_157 ();
 FILLCELL_X2 FILLER_23_166 ();
 FILLCELL_X4 FILLER_23_177 ();
 FILLCELL_X2 FILLER_23_197 ();
 FILLCELL_X1 FILLER_23_199 ();
 FILLCELL_X8 FILLER_23_208 ();
 FILLCELL_X2 FILLER_23_216 ();
 FILLCELL_X2 FILLER_23_224 ();
 FILLCELL_X32 FILLER_23_306 ();
 FILLCELL_X8 FILLER_23_338 ();
 FILLCELL_X2 FILLER_23_372 ();
 FILLCELL_X2 FILLER_23_381 ();
 FILLCELL_X2 FILLER_23_393 ();
 FILLCELL_X1 FILLER_23_395 ();
 FILLCELL_X2 FILLER_23_400 ();
 FILLCELL_X1 FILLER_23_402 ();
 FILLCELL_X1 FILLER_23_409 ();
 FILLCELL_X2 FILLER_23_413 ();
 FILLCELL_X1 FILLER_23_415 ();
 FILLCELL_X2 FILLER_23_426 ();
 FILLCELL_X8 FILLER_23_441 ();
 FILLCELL_X1 FILLER_23_449 ();
 FILLCELL_X2 FILLER_23_461 ();
 FILLCELL_X1 FILLER_23_463 ();
 FILLCELL_X2 FILLER_23_470 ();
 FILLCELL_X4 FILLER_23_476 ();
 FILLCELL_X4 FILLER_23_487 ();
 FILLCELL_X4 FILLER_23_496 ();
 FILLCELL_X1 FILLER_23_500 ();
 FILLCELL_X16 FILLER_23_507 ();
 FILLCELL_X8 FILLER_23_523 ();
 FILLCELL_X4 FILLER_23_531 ();
 FILLCELL_X1 FILLER_23_535 ();
 FILLCELL_X8 FILLER_23_543 ();
 FILLCELL_X4 FILLER_23_551 ();
 FILLCELL_X1 FILLER_23_555 ();
 FILLCELL_X1 FILLER_23_586 ();
 FILLCELL_X2 FILLER_23_615 ();
 FILLCELL_X2 FILLER_23_637 ();
 FILLCELL_X8 FILLER_23_642 ();
 FILLCELL_X2 FILLER_23_650 ();
 FILLCELL_X1 FILLER_23_652 ();
 FILLCELL_X4 FILLER_23_658 ();
 FILLCELL_X1 FILLER_23_662 ();
 FILLCELL_X2 FILLER_23_667 ();
 FILLCELL_X8 FILLER_23_682 ();
 FILLCELL_X2 FILLER_23_690 ();
 FILLCELL_X1 FILLER_23_692 ();
 FILLCELL_X8 FILLER_23_697 ();
 FILLCELL_X2 FILLER_23_705 ();
 FILLCELL_X2 FILLER_23_710 ();
 FILLCELL_X2 FILLER_23_717 ();
 FILLCELL_X2 FILLER_23_723 ();
 FILLCELL_X1 FILLER_23_725 ();
 FILLCELL_X1 FILLER_23_738 ();
 FILLCELL_X4 FILLER_23_745 ();
 FILLCELL_X2 FILLER_23_749 ();
 FILLCELL_X16 FILLER_23_761 ();
 FILLCELL_X8 FILLER_23_777 ();
 FILLCELL_X4 FILLER_23_785 ();
 FILLCELL_X2 FILLER_23_799 ();
 FILLCELL_X2 FILLER_23_817 ();
 FILLCELL_X2 FILLER_23_822 ();
 FILLCELL_X16 FILLER_23_846 ();
 FILLCELL_X4 FILLER_23_866 ();
 FILLCELL_X1 FILLER_23_877 ();
 FILLCELL_X16 FILLER_23_885 ();
 FILLCELL_X4 FILLER_23_901 ();
 FILLCELL_X2 FILLER_23_905 ();
 FILLCELL_X1 FILLER_23_907 ();
 FILLCELL_X4 FILLER_23_915 ();
 FILLCELL_X2 FILLER_23_919 ();
 FILLCELL_X1 FILLER_23_921 ();
 FILLCELL_X2 FILLER_23_943 ();
 FILLCELL_X1 FILLER_23_951 ();
 FILLCELL_X1 FILLER_23_992 ();
 FILLCELL_X1 FILLER_23_1025 ();
 FILLCELL_X4 FILLER_23_1033 ();
 FILLCELL_X2 FILLER_23_1037 ();
 FILLCELL_X1 FILLER_23_1039 ();
 FILLCELL_X32 FILLER_23_1055 ();
 FILLCELL_X32 FILLER_23_1087 ();
 FILLCELL_X32 FILLER_23_1119 ();
 FILLCELL_X32 FILLER_23_1151 ();
 FILLCELL_X16 FILLER_23_1183 ();
 FILLCELL_X8 FILLER_23_1199 ();
 FILLCELL_X2 FILLER_23_1207 ();
 FILLCELL_X32 FILLER_24_1 ();
 FILLCELL_X32 FILLER_24_33 ();
 FILLCELL_X32 FILLER_24_65 ();
 FILLCELL_X32 FILLER_24_97 ();
 FILLCELL_X4 FILLER_24_136 ();
 FILLCELL_X1 FILLER_24_140 ();
 FILLCELL_X1 FILLER_24_164 ();
 FILLCELL_X2 FILLER_24_170 ();
 FILLCELL_X1 FILLER_24_172 ();
 FILLCELL_X1 FILLER_24_177 ();
 FILLCELL_X4 FILLER_24_189 ();
 FILLCELL_X1 FILLER_24_193 ();
 FILLCELL_X2 FILLER_24_200 ();
 FILLCELL_X1 FILLER_24_202 ();
 FILLCELL_X2 FILLER_24_231 ();
 FILLCELL_X2 FILLER_24_247 ();
 FILLCELL_X2 FILLER_24_254 ();
 FILLCELL_X1 FILLER_24_267 ();
 FILLCELL_X2 FILLER_24_286 ();
 FILLCELL_X1 FILLER_24_288 ();
 FILLCELL_X32 FILLER_24_312 ();
 FILLCELL_X4 FILLER_24_344 ();
 FILLCELL_X2 FILLER_24_348 ();
 FILLCELL_X2 FILLER_24_362 ();
 FILLCELL_X1 FILLER_24_364 ();
 FILLCELL_X2 FILLER_24_369 ();
 FILLCELL_X1 FILLER_24_388 ();
 FILLCELL_X8 FILLER_24_402 ();
 FILLCELL_X4 FILLER_24_410 ();
 FILLCELL_X2 FILLER_24_419 ();
 FILLCELL_X2 FILLER_24_429 ();
 FILLCELL_X1 FILLER_24_431 ();
 FILLCELL_X2 FILLER_24_435 ();
 FILLCELL_X1 FILLER_24_437 ();
 FILLCELL_X8 FILLER_24_441 ();
 FILLCELL_X4 FILLER_24_449 ();
 FILLCELL_X2 FILLER_24_453 ();
 FILLCELL_X2 FILLER_24_460 ();
 FILLCELL_X1 FILLER_24_462 ();
 FILLCELL_X2 FILLER_24_467 ();
 FILLCELL_X1 FILLER_24_469 ();
 FILLCELL_X2 FILLER_24_477 ();
 FILLCELL_X1 FILLER_24_490 ();
 FILLCELL_X1 FILLER_24_508 ();
 FILLCELL_X4 FILLER_24_516 ();
 FILLCELL_X1 FILLER_24_520 ();
 FILLCELL_X16 FILLER_24_540 ();
 FILLCELL_X8 FILLER_24_556 ();
 FILLCELL_X1 FILLER_24_564 ();
 FILLCELL_X1 FILLER_24_612 ();
 FILLCELL_X2 FILLER_24_656 ();
 FILLCELL_X4 FILLER_24_672 ();
 FILLCELL_X2 FILLER_24_676 ();
 FILLCELL_X1 FILLER_24_678 ();
 FILLCELL_X2 FILLER_24_701 ();
 FILLCELL_X1 FILLER_24_703 ();
 FILLCELL_X4 FILLER_24_709 ();
 FILLCELL_X2 FILLER_24_713 ();
 FILLCELL_X2 FILLER_24_724 ();
 FILLCELL_X1 FILLER_24_726 ();
 FILLCELL_X2 FILLER_24_735 ();
 FILLCELL_X1 FILLER_24_737 ();
 FILLCELL_X32 FILLER_24_757 ();
 FILLCELL_X8 FILLER_24_789 ();
 FILLCELL_X1 FILLER_24_797 ();
 FILLCELL_X2 FILLER_24_807 ();
 FILLCELL_X2 FILLER_24_848 ();
 FILLCELL_X2 FILLER_24_853 ();
 FILLCELL_X4 FILLER_24_881 ();
 FILLCELL_X32 FILLER_24_895 ();
 FILLCELL_X8 FILLER_24_927 ();
 FILLCELL_X4 FILLER_24_935 ();
 FILLCELL_X2 FILLER_24_939 ();
 FILLCELL_X1 FILLER_24_941 ();
 FILLCELL_X32 FILLER_24_1027 ();
 FILLCELL_X32 FILLER_24_1059 ();
 FILLCELL_X32 FILLER_24_1091 ();
 FILLCELL_X32 FILLER_24_1123 ();
 FILLCELL_X32 FILLER_24_1155 ();
 FILLCELL_X16 FILLER_24_1187 ();
 FILLCELL_X4 FILLER_24_1203 ();
 FILLCELL_X2 FILLER_24_1207 ();
 FILLCELL_X32 FILLER_25_1 ();
 FILLCELL_X32 FILLER_25_33 ();
 FILLCELL_X32 FILLER_25_65 ();
 FILLCELL_X32 FILLER_25_97 ();
 FILLCELL_X1 FILLER_25_129 ();
 FILLCELL_X1 FILLER_25_149 ();
 FILLCELL_X1 FILLER_25_161 ();
 FILLCELL_X1 FILLER_25_165 ();
 FILLCELL_X1 FILLER_25_171 ();
 FILLCELL_X4 FILLER_25_190 ();
 FILLCELL_X2 FILLER_25_194 ();
 FILLCELL_X1 FILLER_25_196 ();
 FILLCELL_X16 FILLER_25_201 ();
 FILLCELL_X4 FILLER_25_217 ();
 FILLCELL_X2 FILLER_25_221 ();
 FILLCELL_X1 FILLER_25_264 ();
 FILLCELL_X4 FILLER_25_304 ();
 FILLCELL_X2 FILLER_25_308 ();
 FILLCELL_X1 FILLER_25_310 ();
 FILLCELL_X8 FILLER_25_336 ();
 FILLCELL_X4 FILLER_25_344 ();
 FILLCELL_X1 FILLER_25_348 ();
 FILLCELL_X8 FILLER_25_365 ();
 FILLCELL_X1 FILLER_25_377 ();
 FILLCELL_X1 FILLER_25_385 ();
 FILLCELL_X2 FILLER_25_398 ();
 FILLCELL_X1 FILLER_25_400 ();
 FILLCELL_X8 FILLER_25_411 ();
 FILLCELL_X1 FILLER_25_419 ();
 FILLCELL_X4 FILLER_25_424 ();
 FILLCELL_X1 FILLER_25_428 ();
 FILLCELL_X4 FILLER_25_436 ();
 FILLCELL_X1 FILLER_25_458 ();
 FILLCELL_X2 FILLER_25_467 ();
 FILLCELL_X1 FILLER_25_473 ();
 FILLCELL_X1 FILLER_25_481 ();
 FILLCELL_X1 FILLER_25_490 ();
 FILLCELL_X16 FILLER_25_505 ();
 FILLCELL_X4 FILLER_25_521 ();
 FILLCELL_X2 FILLER_25_525 ();
 FILLCELL_X1 FILLER_25_527 ();
 FILLCELL_X16 FILLER_25_535 ();
 FILLCELL_X1 FILLER_25_551 ();
 FILLCELL_X4 FILLER_25_560 ();
 FILLCELL_X4 FILLER_25_574 ();
 FILLCELL_X1 FILLER_25_578 ();
 FILLCELL_X2 FILLER_25_620 ();
 FILLCELL_X2 FILLER_25_646 ();
 FILLCELL_X8 FILLER_25_667 ();
 FILLCELL_X4 FILLER_25_675 ();
 FILLCELL_X1 FILLER_25_679 ();
 FILLCELL_X1 FILLER_25_690 ();
 FILLCELL_X2 FILLER_25_701 ();
 FILLCELL_X2 FILLER_25_710 ();
 FILLCELL_X1 FILLER_25_712 ();
 FILLCELL_X4 FILLER_25_716 ();
 FILLCELL_X2 FILLER_25_720 ();
 FILLCELL_X4 FILLER_25_726 ();
 FILLCELL_X1 FILLER_25_730 ();
 FILLCELL_X1 FILLER_25_745 ();
 FILLCELL_X16 FILLER_25_760 ();
 FILLCELL_X8 FILLER_25_776 ();
 FILLCELL_X1 FILLER_25_784 ();
 FILLCELL_X4 FILLER_25_871 ();
 FILLCELL_X2 FILLER_25_897 ();
 FILLCELL_X2 FILLER_25_908 ();
 FILLCELL_X1 FILLER_25_910 ();
 FILLCELL_X1 FILLER_25_915 ();
 FILLCELL_X16 FILLER_25_930 ();
 FILLCELL_X1 FILLER_25_946 ();
 FILLCELL_X1 FILLER_25_954 ();
 FILLCELL_X1 FILLER_25_977 ();
 FILLCELL_X2 FILLER_25_988 ();
 FILLCELL_X32 FILLER_25_1029 ();
 FILLCELL_X32 FILLER_25_1061 ();
 FILLCELL_X32 FILLER_25_1093 ();
 FILLCELL_X32 FILLER_25_1125 ();
 FILLCELL_X32 FILLER_25_1157 ();
 FILLCELL_X16 FILLER_25_1189 ();
 FILLCELL_X4 FILLER_25_1205 ();
 FILLCELL_X32 FILLER_26_1 ();
 FILLCELL_X32 FILLER_26_33 ();
 FILLCELL_X32 FILLER_26_65 ();
 FILLCELL_X16 FILLER_26_97 ();
 FILLCELL_X8 FILLER_26_113 ();
 FILLCELL_X4 FILLER_26_138 ();
 FILLCELL_X1 FILLER_26_149 ();
 FILLCELL_X2 FILLER_26_173 ();
 FILLCELL_X4 FILLER_26_179 ();
 FILLCELL_X2 FILLER_26_183 ();
 FILLCELL_X2 FILLER_26_188 ();
 FILLCELL_X1 FILLER_26_190 ();
 FILLCELL_X2 FILLER_26_200 ();
 FILLCELL_X1 FILLER_26_202 ();
 FILLCELL_X8 FILLER_26_206 ();
 FILLCELL_X4 FILLER_26_214 ();
 FILLCELL_X1 FILLER_26_218 ();
 FILLCELL_X2 FILLER_26_246 ();
 FILLCELL_X2 FILLER_26_252 ();
 FILLCELL_X1 FILLER_26_262 ();
 FILLCELL_X2 FILLER_26_266 ();
 FILLCELL_X1 FILLER_26_286 ();
 FILLCELL_X32 FILLER_26_308 ();
 FILLCELL_X8 FILLER_26_340 ();
 FILLCELL_X2 FILLER_26_355 ();
 FILLCELL_X2 FILLER_26_373 ();
 FILLCELL_X1 FILLER_26_375 ();
 FILLCELL_X8 FILLER_26_395 ();
 FILLCELL_X1 FILLER_26_403 ();
 FILLCELL_X4 FILLER_26_408 ();
 FILLCELL_X1 FILLER_26_412 ();
 FILLCELL_X4 FILLER_26_418 ();
 FILLCELL_X1 FILLER_26_422 ();
 FILLCELL_X8 FILLER_26_427 ();
 FILLCELL_X4 FILLER_26_435 ();
 FILLCELL_X1 FILLER_26_439 ();
 FILLCELL_X1 FILLER_26_447 ();
 FILLCELL_X1 FILLER_26_463 ();
 FILLCELL_X2 FILLER_26_497 ();
 FILLCELL_X1 FILLER_26_499 ();
 FILLCELL_X16 FILLER_26_504 ();
 FILLCELL_X4 FILLER_26_520 ();
 FILLCELL_X2 FILLER_26_524 ();
 FILLCELL_X16 FILLER_26_543 ();
 FILLCELL_X8 FILLER_26_559 ();
 FILLCELL_X1 FILLER_26_567 ();
 FILLCELL_X1 FILLER_26_604 ();
 FILLCELL_X2 FILLER_26_612 ();
 FILLCELL_X2 FILLER_26_628 ();
 FILLCELL_X1 FILLER_26_630 ();
 FILLCELL_X8 FILLER_26_632 ();
 FILLCELL_X1 FILLER_26_640 ();
 FILLCELL_X2 FILLER_26_648 ();
 FILLCELL_X1 FILLER_26_650 ();
 FILLCELL_X1 FILLER_26_654 ();
 FILLCELL_X2 FILLER_26_658 ();
 FILLCELL_X1 FILLER_26_660 ();
 FILLCELL_X4 FILLER_26_664 ();
 FILLCELL_X2 FILLER_26_668 ();
 FILLCELL_X8 FILLER_26_674 ();
 FILLCELL_X4 FILLER_26_682 ();
 FILLCELL_X8 FILLER_26_696 ();
 FILLCELL_X1 FILLER_26_704 ();
 FILLCELL_X2 FILLER_26_717 ();
 FILLCELL_X2 FILLER_26_727 ();
 FILLCELL_X4 FILLER_26_745 ();
 FILLCELL_X2 FILLER_26_749 ();
 FILLCELL_X16 FILLER_26_755 ();
 FILLCELL_X4 FILLER_26_771 ();
 FILLCELL_X2 FILLER_26_775 ();
 FILLCELL_X4 FILLER_26_787 ();
 FILLCELL_X2 FILLER_26_791 ();
 FILLCELL_X1 FILLER_26_793 ();
 FILLCELL_X1 FILLER_26_884 ();
 FILLCELL_X2 FILLER_26_893 ();
 FILLCELL_X1 FILLER_26_895 ();
 FILLCELL_X4 FILLER_26_901 ();
 FILLCELL_X2 FILLER_26_905 ();
 FILLCELL_X16 FILLER_26_929 ();
 FILLCELL_X8 FILLER_26_945 ();
 FILLCELL_X2 FILLER_26_956 ();
 FILLCELL_X2 FILLER_26_961 ();
 FILLCELL_X1 FILLER_26_963 ();
 FILLCELL_X2 FILLER_26_974 ();
 FILLCELL_X32 FILLER_26_1024 ();
 FILLCELL_X32 FILLER_26_1056 ();
 FILLCELL_X32 FILLER_26_1088 ();
 FILLCELL_X32 FILLER_26_1120 ();
 FILLCELL_X32 FILLER_26_1152 ();
 FILLCELL_X16 FILLER_26_1184 ();
 FILLCELL_X8 FILLER_26_1200 ();
 FILLCELL_X1 FILLER_26_1208 ();
 FILLCELL_X32 FILLER_27_1 ();
 FILLCELL_X32 FILLER_27_33 ();
 FILLCELL_X32 FILLER_27_65 ();
 FILLCELL_X32 FILLER_27_97 ();
 FILLCELL_X2 FILLER_27_129 ();
 FILLCELL_X2 FILLER_27_136 ();
 FILLCELL_X1 FILLER_27_138 ();
 FILLCELL_X2 FILLER_27_169 ();
 FILLCELL_X1 FILLER_27_171 ();
 FILLCELL_X4 FILLER_27_175 ();
 FILLCELL_X2 FILLER_27_190 ();
 FILLCELL_X1 FILLER_27_201 ();
 FILLCELL_X1 FILLER_27_227 ();
 FILLCELL_X2 FILLER_27_235 ();
 FILLCELL_X8 FILLER_27_250 ();
 FILLCELL_X4 FILLER_27_258 ();
 FILLCELL_X2 FILLER_27_262 ();
 FILLCELL_X32 FILLER_27_318 ();
 FILLCELL_X8 FILLER_27_350 ();
 FILLCELL_X4 FILLER_27_358 ();
 FILLCELL_X1 FILLER_27_362 ();
 FILLCELL_X1 FILLER_27_375 ();
 FILLCELL_X4 FILLER_27_405 ();
 FILLCELL_X2 FILLER_27_421 ();
 FILLCELL_X1 FILLER_27_423 ();
 FILLCELL_X1 FILLER_27_428 ();
 FILLCELL_X2 FILLER_27_451 ();
 FILLCELL_X1 FILLER_27_453 ();
 FILLCELL_X8 FILLER_27_460 ();
 FILLCELL_X2 FILLER_27_468 ();
 FILLCELL_X1 FILLER_27_470 ();
 FILLCELL_X2 FILLER_27_475 ();
 FILLCELL_X1 FILLER_27_483 ();
 FILLCELL_X32 FILLER_27_498 ();
 FILLCELL_X1 FILLER_27_530 ();
 FILLCELL_X32 FILLER_27_538 ();
 FILLCELL_X2 FILLER_27_582 ();
 FILLCELL_X1 FILLER_27_611 ();
 FILLCELL_X8 FILLER_27_669 ();
 FILLCELL_X1 FILLER_27_691 ();
 FILLCELL_X8 FILLER_27_699 ();
 FILLCELL_X1 FILLER_27_707 ();
 FILLCELL_X8 FILLER_27_711 ();
 FILLCELL_X4 FILLER_27_719 ();
 FILLCELL_X2 FILLER_27_723 ();
 FILLCELL_X1 FILLER_27_733 ();
 FILLCELL_X4 FILLER_27_748 ();
 FILLCELL_X2 FILLER_27_752 ();
 FILLCELL_X32 FILLER_27_764 ();
 FILLCELL_X8 FILLER_27_796 ();
 FILLCELL_X2 FILLER_27_804 ();
 FILLCELL_X1 FILLER_27_806 ();
 FILLCELL_X1 FILLER_27_845 ();
 FILLCELL_X2 FILLER_27_853 ();
 FILLCELL_X1 FILLER_27_877 ();
 FILLCELL_X1 FILLER_27_896 ();
 FILLCELL_X1 FILLER_27_918 ();
 FILLCELL_X16 FILLER_27_938 ();
 FILLCELL_X8 FILLER_27_954 ();
 FILLCELL_X4 FILLER_27_962 ();
 FILLCELL_X2 FILLER_27_966 ();
 FILLCELL_X1 FILLER_27_968 ();
 FILLCELL_X2 FILLER_27_998 ();
 FILLCELL_X32 FILLER_27_1017 ();
 FILLCELL_X32 FILLER_27_1049 ();
 FILLCELL_X32 FILLER_27_1081 ();
 FILLCELL_X32 FILLER_27_1113 ();
 FILLCELL_X32 FILLER_27_1145 ();
 FILLCELL_X32 FILLER_27_1177 ();
 FILLCELL_X32 FILLER_28_1 ();
 FILLCELL_X32 FILLER_28_33 ();
 FILLCELL_X32 FILLER_28_65 ();
 FILLCELL_X32 FILLER_28_97 ();
 FILLCELL_X2 FILLER_28_129 ();
 FILLCELL_X1 FILLER_28_131 ();
 FILLCELL_X2 FILLER_28_168 ();
 FILLCELL_X2 FILLER_28_191 ();
 FILLCELL_X1 FILLER_28_196 ();
 FILLCELL_X2 FILLER_28_202 ();
 FILLCELL_X1 FILLER_28_204 ();
 FILLCELL_X4 FILLER_28_237 ();
 FILLCELL_X2 FILLER_28_241 ();
 FILLCELL_X1 FILLER_28_243 ();
 FILLCELL_X1 FILLER_28_251 ();
 FILLCELL_X4 FILLER_28_256 ();
 FILLCELL_X4 FILLER_28_266 ();
 FILLCELL_X1 FILLER_28_270 ();
 FILLCELL_X2 FILLER_28_286 ();
 FILLCELL_X32 FILLER_28_314 ();
 FILLCELL_X4 FILLER_28_354 ();
 FILLCELL_X1 FILLER_28_358 ();
 FILLCELL_X2 FILLER_28_364 ();
 FILLCELL_X4 FILLER_28_389 ();
 FILLCELL_X8 FILLER_28_420 ();
 FILLCELL_X8 FILLER_28_434 ();
 FILLCELL_X4 FILLER_28_447 ();
 FILLCELL_X2 FILLER_28_451 ();
 FILLCELL_X1 FILLER_28_479 ();
 FILLCELL_X2 FILLER_28_498 ();
 FILLCELL_X8 FILLER_28_505 ();
 FILLCELL_X2 FILLER_28_513 ();
 FILLCELL_X1 FILLER_28_515 ();
 FILLCELL_X16 FILLER_28_533 ();
 FILLCELL_X4 FILLER_28_549 ();
 FILLCELL_X1 FILLER_28_553 ();
 FILLCELL_X1 FILLER_28_573 ();
 FILLCELL_X4 FILLER_28_623 ();
 FILLCELL_X2 FILLER_28_641 ();
 FILLCELL_X1 FILLER_28_643 ();
 FILLCELL_X8 FILLER_28_668 ();
 FILLCELL_X1 FILLER_28_676 ();
 FILLCELL_X1 FILLER_28_705 ();
 FILLCELL_X1 FILLER_28_713 ();
 FILLCELL_X4 FILLER_28_730 ();
 FILLCELL_X32 FILLER_28_738 ();
 FILLCELL_X8 FILLER_28_770 ();
 FILLCELL_X4 FILLER_28_783 ();
 FILLCELL_X2 FILLER_28_787 ();
 FILLCELL_X1 FILLER_28_799 ();
 FILLCELL_X2 FILLER_28_816 ();
 FILLCELL_X2 FILLER_28_842 ();
 FILLCELL_X1 FILLER_28_844 ();
 FILLCELL_X4 FILLER_28_870 ();
 FILLCELL_X2 FILLER_28_890 ();
 FILLCELL_X1 FILLER_28_901 ();
 FILLCELL_X2 FILLER_28_915 ();
 FILLCELL_X4 FILLER_28_924 ();
 FILLCELL_X16 FILLER_28_938 ();
 FILLCELL_X8 FILLER_28_954 ();
 FILLCELL_X4 FILLER_28_962 ();
 FILLCELL_X2 FILLER_28_966 ();
 FILLCELL_X1 FILLER_28_968 ();
 FILLCELL_X1 FILLER_28_987 ();
 FILLCELL_X2 FILLER_28_991 ();
 FILLCELL_X1 FILLER_28_993 ();
 FILLCELL_X2 FILLER_28_997 ();
 FILLCELL_X32 FILLER_28_1018 ();
 FILLCELL_X16 FILLER_28_1050 ();
 FILLCELL_X4 FILLER_28_1066 ();
 FILLCELL_X2 FILLER_28_1070 ();
 FILLCELL_X32 FILLER_28_1079 ();
 FILLCELL_X8 FILLER_28_1111 ();
 FILLCELL_X2 FILLER_28_1119 ();
 FILLCELL_X1 FILLER_28_1121 ();
 FILLCELL_X32 FILLER_28_1171 ();
 FILLCELL_X4 FILLER_28_1203 ();
 FILLCELL_X2 FILLER_28_1207 ();
 FILLCELL_X32 FILLER_29_1 ();
 FILLCELL_X32 FILLER_29_33 ();
 FILLCELL_X32 FILLER_29_65 ();
 FILLCELL_X32 FILLER_29_97 ();
 FILLCELL_X16 FILLER_29_129 ();
 FILLCELL_X2 FILLER_29_145 ();
 FILLCELL_X4 FILLER_29_151 ();
 FILLCELL_X2 FILLER_29_164 ();
 FILLCELL_X1 FILLER_29_166 ();
 FILLCELL_X2 FILLER_29_184 ();
 FILLCELL_X4 FILLER_29_204 ();
 FILLCELL_X1 FILLER_29_218 ();
 FILLCELL_X8 FILLER_29_226 ();
 FILLCELL_X1 FILLER_29_234 ();
 FILLCELL_X1 FILLER_29_267 ();
 FILLCELL_X2 FILLER_29_278 ();
 FILLCELL_X1 FILLER_29_280 ();
 FILLCELL_X2 FILLER_29_292 ();
 FILLCELL_X32 FILLER_29_308 ();
 FILLCELL_X4 FILLER_29_340 ();
 FILLCELL_X2 FILLER_29_344 ();
 FILLCELL_X1 FILLER_29_346 ();
 FILLCELL_X2 FILLER_29_356 ();
 FILLCELL_X1 FILLER_29_358 ();
 FILLCELL_X1 FILLER_29_368 ();
 FILLCELL_X1 FILLER_29_373 ();
 FILLCELL_X1 FILLER_29_382 ();
 FILLCELL_X2 FILLER_29_394 ();
 FILLCELL_X2 FILLER_29_405 ();
 FILLCELL_X4 FILLER_29_419 ();
 FILLCELL_X2 FILLER_29_430 ();
 FILLCELL_X1 FILLER_29_450 ();
 FILLCELL_X4 FILLER_29_466 ();
 FILLCELL_X1 FILLER_29_470 ();
 FILLCELL_X2 FILLER_29_474 ();
 FILLCELL_X1 FILLER_29_480 ();
 FILLCELL_X16 FILLER_29_499 ();
 FILLCELL_X4 FILLER_29_515 ();
 FILLCELL_X4 FILLER_29_568 ();
 FILLCELL_X1 FILLER_29_572 ();
 FILLCELL_X16 FILLER_29_596 ();
 FILLCELL_X4 FILLER_29_612 ();
 FILLCELL_X2 FILLER_29_616 ();
 FILLCELL_X1 FILLER_29_618 ();
 FILLCELL_X1 FILLER_29_629 ();
 FILLCELL_X1 FILLER_29_666 ();
 FILLCELL_X8 FILLER_29_672 ();
 FILLCELL_X2 FILLER_29_690 ();
 FILLCELL_X32 FILLER_29_722 ();
 FILLCELL_X8 FILLER_29_754 ();
 FILLCELL_X2 FILLER_29_762 ();
 FILLCELL_X1 FILLER_29_764 ();
 FILLCELL_X4 FILLER_29_785 ();
 FILLCELL_X2 FILLER_29_789 ();
 FILLCELL_X1 FILLER_29_802 ();
 FILLCELL_X2 FILLER_29_808 ();
 FILLCELL_X1 FILLER_29_810 ();
 FILLCELL_X2 FILLER_29_836 ();
 FILLCELL_X1 FILLER_29_838 ();
 FILLCELL_X1 FILLER_29_850 ();
 FILLCELL_X2 FILLER_29_876 ();
 FILLCELL_X1 FILLER_29_878 ();
 FILLCELL_X2 FILLER_29_893 ();
 FILLCELL_X1 FILLER_29_905 ();
 FILLCELL_X2 FILLER_29_920 ();
 FILLCELL_X8 FILLER_29_941 ();
 FILLCELL_X4 FILLER_29_949 ();
 FILLCELL_X2 FILLER_29_953 ();
 FILLCELL_X2 FILLER_29_964 ();
 FILLCELL_X1 FILLER_29_966 ();
 FILLCELL_X32 FILLER_29_999 ();
 FILLCELL_X1 FILLER_29_1031 ();
 FILLCELL_X4 FILLER_29_1082 ();
 FILLCELL_X1 FILLER_29_1086 ();
 FILLCELL_X32 FILLER_29_1112 ();
 FILLCELL_X32 FILLER_29_1144 ();
 FILLCELL_X32 FILLER_29_1176 ();
 FILLCELL_X1 FILLER_29_1208 ();
 FILLCELL_X32 FILLER_30_1 ();
 FILLCELL_X32 FILLER_30_33 ();
 FILLCELL_X32 FILLER_30_65 ();
 FILLCELL_X32 FILLER_30_97 ();
 FILLCELL_X8 FILLER_30_129 ();
 FILLCELL_X2 FILLER_30_137 ();
 FILLCELL_X1 FILLER_30_151 ();
 FILLCELL_X2 FILLER_30_161 ();
 FILLCELL_X1 FILLER_30_163 ();
 FILLCELL_X4 FILLER_30_169 ();
 FILLCELL_X16 FILLER_30_185 ();
 FILLCELL_X8 FILLER_30_201 ();
 FILLCELL_X1 FILLER_30_209 ();
 FILLCELL_X4 FILLER_30_220 ();
 FILLCELL_X1 FILLER_30_224 ();
 FILLCELL_X1 FILLER_30_233 ();
 FILLCELL_X1 FILLER_30_238 ();
 FILLCELL_X1 FILLER_30_261 ();
 FILLCELL_X1 FILLER_30_272 ();
 FILLCELL_X8 FILLER_30_280 ();
 FILLCELL_X4 FILLER_30_288 ();
 FILLCELL_X2 FILLER_30_292 ();
 FILLCELL_X16 FILLER_30_301 ();
 FILLCELL_X2 FILLER_30_317 ();
 FILLCELL_X1 FILLER_30_319 ();
 FILLCELL_X4 FILLER_30_330 ();
 FILLCELL_X1 FILLER_30_334 ();
 FILLCELL_X32 FILLER_30_338 ();
 FILLCELL_X2 FILLER_30_370 ();
 FILLCELL_X1 FILLER_30_372 ();
 FILLCELL_X4 FILLER_30_380 ();
 FILLCELL_X2 FILLER_30_384 ();
 FILLCELL_X1 FILLER_30_386 ();
 FILLCELL_X4 FILLER_30_396 ();
 FILLCELL_X1 FILLER_30_400 ();
 FILLCELL_X1 FILLER_30_410 ();
 FILLCELL_X4 FILLER_30_432 ();
 FILLCELL_X4 FILLER_30_439 ();
 FILLCELL_X1 FILLER_30_443 ();
 FILLCELL_X4 FILLER_30_462 ();
 FILLCELL_X1 FILLER_30_469 ();
 FILLCELL_X2 FILLER_30_475 ();
 FILLCELL_X2 FILLER_30_486 ();
 FILLCELL_X32 FILLER_30_502 ();
 FILLCELL_X4 FILLER_30_534 ();
 FILLCELL_X2 FILLER_30_538 ();
 FILLCELL_X2 FILLER_30_553 ();
 FILLCELL_X4 FILLER_30_575 ();
 FILLCELL_X2 FILLER_30_579 ();
 FILLCELL_X1 FILLER_30_581 ();
 FILLCELL_X2 FILLER_30_605 ();
 FILLCELL_X1 FILLER_30_607 ();
 FILLCELL_X1 FILLER_30_648 ();
 FILLCELL_X1 FILLER_30_658 ();
 FILLCELL_X4 FILLER_30_674 ();
 FILLCELL_X2 FILLER_30_678 ();
 FILLCELL_X1 FILLER_30_680 ();
 FILLCELL_X2 FILLER_30_695 ();
 FILLCELL_X8 FILLER_30_703 ();
 FILLCELL_X4 FILLER_30_711 ();
 FILLCELL_X2 FILLER_30_715 ();
 FILLCELL_X1 FILLER_30_717 ();
 FILLCELL_X4 FILLER_30_722 ();
 FILLCELL_X2 FILLER_30_726 ();
 FILLCELL_X1 FILLER_30_728 ();
 FILLCELL_X16 FILLER_30_743 ();
 FILLCELL_X8 FILLER_30_784 ();
 FILLCELL_X4 FILLER_30_797 ();
 FILLCELL_X2 FILLER_30_801 ();
 FILLCELL_X2 FILLER_30_859 ();
 FILLCELL_X1 FILLER_30_861 ();
 FILLCELL_X1 FILLER_30_882 ();
 FILLCELL_X2 FILLER_30_928 ();
 FILLCELL_X8 FILLER_30_943 ();
 FILLCELL_X4 FILLER_30_951 ();
 FILLCELL_X1 FILLER_30_955 ();
 FILLCELL_X2 FILLER_30_966 ();
 FILLCELL_X1 FILLER_30_968 ();
 FILLCELL_X32 FILLER_30_983 ();
 FILLCELL_X16 FILLER_30_1015 ();
 FILLCELL_X1 FILLER_30_1031 ();
 FILLCELL_X8 FILLER_30_1058 ();
 FILLCELL_X8 FILLER_30_1118 ();
 FILLCELL_X2 FILLER_30_1133 ();
 FILLCELL_X1 FILLER_30_1135 ();
 FILLCELL_X4 FILLER_30_1143 ();
 FILLCELL_X1 FILLER_30_1147 ();
 FILLCELL_X32 FILLER_30_1173 ();
 FILLCELL_X4 FILLER_30_1205 ();
 FILLCELL_X32 FILLER_31_1 ();
 FILLCELL_X32 FILLER_31_33 ();
 FILLCELL_X32 FILLER_31_65 ();
 FILLCELL_X32 FILLER_31_97 ();
 FILLCELL_X8 FILLER_31_129 ();
 FILLCELL_X2 FILLER_31_137 ();
 FILLCELL_X1 FILLER_31_139 ();
 FILLCELL_X1 FILLER_31_147 ();
 FILLCELL_X1 FILLER_31_171 ();
 FILLCELL_X1 FILLER_31_179 ();
 FILLCELL_X4 FILLER_31_194 ();
 FILLCELL_X2 FILLER_31_198 ();
 FILLCELL_X1 FILLER_31_200 ();
 FILLCELL_X8 FILLER_31_205 ();
 FILLCELL_X1 FILLER_31_213 ();
 FILLCELL_X4 FILLER_31_219 ();
 FILLCELL_X4 FILLER_31_232 ();
 FILLCELL_X1 FILLER_31_236 ();
 FILLCELL_X2 FILLER_31_241 ();
 FILLCELL_X1 FILLER_31_250 ();
 FILLCELL_X1 FILLER_31_254 ();
 FILLCELL_X2 FILLER_31_260 ();
 FILLCELL_X8 FILLER_31_267 ();
 FILLCELL_X4 FILLER_31_275 ();
 FILLCELL_X16 FILLER_31_300 ();
 FILLCELL_X4 FILLER_31_316 ();
 FILLCELL_X2 FILLER_31_320 ();
 FILLCELL_X32 FILLER_31_355 ();
 FILLCELL_X2 FILLER_31_387 ();
 FILLCELL_X4 FILLER_31_396 ();
 FILLCELL_X2 FILLER_31_400 ();
 FILLCELL_X16 FILLER_31_407 ();
 FILLCELL_X8 FILLER_31_423 ();
 FILLCELL_X1 FILLER_31_431 ();
 FILLCELL_X8 FILLER_31_436 ();
 FILLCELL_X4 FILLER_31_453 ();
 FILLCELL_X2 FILLER_31_457 ();
 FILLCELL_X2 FILLER_31_473 ();
 FILLCELL_X2 FILLER_31_478 ();
 FILLCELL_X32 FILLER_31_487 ();
 FILLCELL_X32 FILLER_31_519 ();
 FILLCELL_X4 FILLER_31_551 ();
 FILLCELL_X8 FILLER_31_568 ();
 FILLCELL_X1 FILLER_31_576 ();
 FILLCELL_X2 FILLER_31_598 ();
 FILLCELL_X1 FILLER_31_600 ();
 FILLCELL_X4 FILLER_31_614 ();
 FILLCELL_X2 FILLER_31_618 ();
 FILLCELL_X1 FILLER_31_620 ();
 FILLCELL_X4 FILLER_31_651 ();
 FILLCELL_X2 FILLER_31_655 ();
 FILLCELL_X16 FILLER_31_663 ();
 FILLCELL_X4 FILLER_31_679 ();
 FILLCELL_X2 FILLER_31_683 ();
 FILLCELL_X1 FILLER_31_685 ();
 FILLCELL_X1 FILLER_31_697 ();
 FILLCELL_X1 FILLER_31_702 ();
 FILLCELL_X4 FILLER_31_711 ();
 FILLCELL_X1 FILLER_31_715 ();
 FILLCELL_X2 FILLER_31_721 ();
 FILLCELL_X16 FILLER_31_729 ();
 FILLCELL_X8 FILLER_31_745 ();
 FILLCELL_X2 FILLER_31_863 ();
 FILLCELL_X1 FILLER_31_865 ();
 FILLCELL_X1 FILLER_31_871 ();
 FILLCELL_X1 FILLER_31_895 ();
 FILLCELL_X1 FILLER_31_900 ();
 FILLCELL_X1 FILLER_31_909 ();
 FILLCELL_X8 FILLER_31_947 ();
 FILLCELL_X2 FILLER_31_955 ();
 FILLCELL_X1 FILLER_31_957 ();
 FILLCELL_X8 FILLER_31_967 ();
 FILLCELL_X4 FILLER_31_975 ();
 FILLCELL_X2 FILLER_31_979 ();
 FILLCELL_X16 FILLER_31_1000 ();
 FILLCELL_X8 FILLER_31_1016 ();
 FILLCELL_X2 FILLER_31_1024 ();
 FILLCELL_X1 FILLER_31_1026 ();
 FILLCELL_X4 FILLER_31_1048 ();
 FILLCELL_X4 FILLER_31_1059 ();
 FILLCELL_X1 FILLER_31_1063 ();
 FILLCELL_X4 FILLER_31_1074 ();
 FILLCELL_X1 FILLER_31_1078 ();
 FILLCELL_X1 FILLER_31_1097 ();
 FILLCELL_X1 FILLER_31_1128 ();
 FILLCELL_X2 FILLER_31_1136 ();
 FILLCELL_X2 FILLER_31_1142 ();
 FILLCELL_X4 FILLER_31_1148 ();
 FILLCELL_X2 FILLER_31_1152 ();
 FILLCELL_X1 FILLER_31_1154 ();
 FILLCELL_X2 FILLER_31_1165 ();
 FILLCELL_X16 FILLER_31_1192 ();
 FILLCELL_X1 FILLER_31_1208 ();
 FILLCELL_X32 FILLER_32_1 ();
 FILLCELL_X32 FILLER_32_33 ();
 FILLCELL_X32 FILLER_32_65 ();
 FILLCELL_X32 FILLER_32_97 ();
 FILLCELL_X16 FILLER_32_129 ();
 FILLCELL_X8 FILLER_32_145 ();
 FILLCELL_X2 FILLER_32_153 ();
 FILLCELL_X1 FILLER_32_155 ();
 FILLCELL_X2 FILLER_32_181 ();
 FILLCELL_X1 FILLER_32_183 ();
 FILLCELL_X1 FILLER_32_186 ();
 FILLCELL_X1 FILLER_32_191 ();
 FILLCELL_X2 FILLER_32_196 ();
 FILLCELL_X1 FILLER_32_202 ();
 FILLCELL_X2 FILLER_32_238 ();
 FILLCELL_X8 FILLER_32_245 ();
 FILLCELL_X2 FILLER_32_253 ();
 FILLCELL_X16 FILLER_32_262 ();
 FILLCELL_X4 FILLER_32_278 ();
 FILLCELL_X16 FILLER_32_301 ();
 FILLCELL_X4 FILLER_32_336 ();
 FILLCELL_X2 FILLER_32_340 ();
 FILLCELL_X1 FILLER_32_342 ();
 FILLCELL_X4 FILLER_32_377 ();
 FILLCELL_X2 FILLER_32_381 ();
 FILLCELL_X1 FILLER_32_383 ();
 FILLCELL_X32 FILLER_32_408 ();
 FILLCELL_X16 FILLER_32_440 ();
 FILLCELL_X1 FILLER_32_456 ();
 FILLCELL_X4 FILLER_32_464 ();
 FILLCELL_X1 FILLER_32_468 ();
 FILLCELL_X8 FILLER_32_488 ();
 FILLCELL_X4 FILLER_32_522 ();
 FILLCELL_X2 FILLER_32_526 ();
 FILLCELL_X16 FILLER_32_537 ();
 FILLCELL_X8 FILLER_32_553 ();
 FILLCELL_X4 FILLER_32_561 ();
 FILLCELL_X2 FILLER_32_565 ();
 FILLCELL_X1 FILLER_32_567 ();
 FILLCELL_X4 FILLER_32_594 ();
 FILLCELL_X1 FILLER_32_598 ();
 FILLCELL_X2 FILLER_32_606 ();
 FILLCELL_X1 FILLER_32_615 ();
 FILLCELL_X2 FILLER_32_620 ();
 FILLCELL_X1 FILLER_32_632 ();
 FILLCELL_X4 FILLER_32_648 ();
 FILLCELL_X2 FILLER_32_652 ();
 FILLCELL_X1 FILLER_32_654 ();
 FILLCELL_X8 FILLER_32_669 ();
 FILLCELL_X4 FILLER_32_677 ();
 FILLCELL_X2 FILLER_32_681 ();
 FILLCELL_X1 FILLER_32_683 ();
 FILLCELL_X16 FILLER_32_691 ();
 FILLCELL_X8 FILLER_32_707 ();
 FILLCELL_X16 FILLER_32_722 ();
 FILLCELL_X8 FILLER_32_738 ();
 FILLCELL_X4 FILLER_32_746 ();
 FILLCELL_X2 FILLER_32_750 ();
 FILLCELL_X4 FILLER_32_781 ();
 FILLCELL_X2 FILLER_32_785 ();
 FILLCELL_X1 FILLER_32_787 ();
 FILLCELL_X2 FILLER_32_827 ();
 FILLCELL_X1 FILLER_32_829 ();
 FILLCELL_X2 FILLER_32_862 ();
 FILLCELL_X4 FILLER_32_876 ();
 FILLCELL_X2 FILLER_32_880 ();
 FILLCELL_X1 FILLER_32_882 ();
 FILLCELL_X4 FILLER_32_946 ();
 FILLCELL_X2 FILLER_32_950 ();
 FILLCELL_X1 FILLER_32_952 ();
 FILLCELL_X16 FILLER_32_974 ();
 FILLCELL_X2 FILLER_32_990 ();
 FILLCELL_X8 FILLER_32_1013 ();
 FILLCELL_X2 FILLER_32_1021 ();
 FILLCELL_X1 FILLER_32_1023 ();
 FILLCELL_X2 FILLER_32_1054 ();
 FILLCELL_X2 FILLER_32_1092 ();
 FILLCELL_X2 FILLER_32_1129 ();
 FILLCELL_X1 FILLER_32_1131 ();
 FILLCELL_X1 FILLER_32_1146 ();
 FILLCELL_X8 FILLER_32_1164 ();
 FILLCELL_X16 FILLER_32_1185 ();
 FILLCELL_X8 FILLER_32_1201 ();
 FILLCELL_X32 FILLER_33_1 ();
 FILLCELL_X32 FILLER_33_33 ();
 FILLCELL_X32 FILLER_33_65 ();
 FILLCELL_X32 FILLER_33_97 ();
 FILLCELL_X16 FILLER_33_129 ();
 FILLCELL_X8 FILLER_33_145 ();
 FILLCELL_X4 FILLER_33_153 ();
 FILLCELL_X1 FILLER_33_157 ();
 FILLCELL_X4 FILLER_33_169 ();
 FILLCELL_X1 FILLER_33_173 ();
 FILLCELL_X2 FILLER_33_192 ();
 FILLCELL_X2 FILLER_33_213 ();
 FILLCELL_X1 FILLER_33_215 ();
 FILLCELL_X1 FILLER_33_227 ();
 FILLCELL_X4 FILLER_33_237 ();
 FILLCELL_X1 FILLER_33_254 ();
 FILLCELL_X2 FILLER_33_260 ();
 FILLCELL_X1 FILLER_33_262 ();
 FILLCELL_X4 FILLER_33_276 ();
 FILLCELL_X1 FILLER_33_280 ();
 FILLCELL_X4 FILLER_33_288 ();
 FILLCELL_X1 FILLER_33_292 ();
 FILLCELL_X2 FILLER_33_302 ();
 FILLCELL_X8 FILLER_33_350 ();
 FILLCELL_X2 FILLER_33_363 ();
 FILLCELL_X16 FILLER_33_371 ();
 FILLCELL_X8 FILLER_33_387 ();
 FILLCELL_X4 FILLER_33_395 ();
 FILLCELL_X1 FILLER_33_399 ();
 FILLCELL_X2 FILLER_33_405 ();
 FILLCELL_X2 FILLER_33_424 ();
 FILLCELL_X4 FILLER_33_443 ();
 FILLCELL_X2 FILLER_33_464 ();
 FILLCELL_X2 FILLER_33_475 ();
 FILLCELL_X4 FILLER_33_482 ();
 FILLCELL_X4 FILLER_33_503 ();
 FILLCELL_X4 FILLER_33_512 ();
 FILLCELL_X16 FILLER_33_532 ();
 FILLCELL_X1 FILLER_33_548 ();
 FILLCELL_X8 FILLER_33_556 ();
 FILLCELL_X4 FILLER_33_564 ();
 FILLCELL_X1 FILLER_33_568 ();
 FILLCELL_X2 FILLER_33_596 ();
 FILLCELL_X4 FILLER_33_611 ();
 FILLCELL_X2 FILLER_33_615 ();
 FILLCELL_X2 FILLER_33_634 ();
 FILLCELL_X1 FILLER_33_636 ();
 FILLCELL_X8 FILLER_33_641 ();
 FILLCELL_X2 FILLER_33_649 ();
 FILLCELL_X4 FILLER_33_661 ();
 FILLCELL_X2 FILLER_33_665 ();
 FILLCELL_X1 FILLER_33_667 ();
 FILLCELL_X1 FILLER_33_675 ();
 FILLCELL_X4 FILLER_33_679 ();
 FILLCELL_X32 FILLER_33_697 ();
 FILLCELL_X16 FILLER_33_729 ();
 FILLCELL_X8 FILLER_33_745 ();
 FILLCELL_X2 FILLER_33_753 ();
 FILLCELL_X2 FILLER_33_788 ();
 FILLCELL_X2 FILLER_33_821 ();
 FILLCELL_X1 FILLER_33_849 ();
 FILLCELL_X2 FILLER_33_862 ();
 FILLCELL_X4 FILLER_33_875 ();
 FILLCELL_X8 FILLER_33_883 ();
 FILLCELL_X4 FILLER_33_891 ();
 FILLCELL_X1 FILLER_33_895 ();
 FILLCELL_X2 FILLER_33_936 ();
 FILLCELL_X8 FILLER_33_943 ();
 FILLCELL_X4 FILLER_33_951 ();
 FILLCELL_X2 FILLER_33_955 ();
 FILLCELL_X4 FILLER_33_973 ();
 FILLCELL_X2 FILLER_33_977 ();
 FILLCELL_X16 FILLER_33_988 ();
 FILLCELL_X4 FILLER_33_1004 ();
 FILLCELL_X2 FILLER_33_1008 ();
 FILLCELL_X16 FILLER_33_1017 ();
 FILLCELL_X4 FILLER_33_1047 ();
 FILLCELL_X2 FILLER_33_1051 ();
 FILLCELL_X2 FILLER_33_1071 ();
 FILLCELL_X2 FILLER_33_1076 ();
 FILLCELL_X1 FILLER_33_1078 ();
 FILLCELL_X1 FILLER_33_1086 ();
 FILLCELL_X2 FILLER_33_1094 ();
 FILLCELL_X1 FILLER_33_1105 ();
 FILLCELL_X2 FILLER_33_1125 ();
 FILLCELL_X1 FILLER_33_1127 ();
 FILLCELL_X2 FILLER_33_1136 ();
 FILLCELL_X2 FILLER_33_1148 ();
 FILLCELL_X1 FILLER_33_1150 ();
 FILLCELL_X1 FILLER_33_1159 ();
 FILLCELL_X2 FILLER_33_1170 ();
 FILLCELL_X32 FILLER_33_1177 ();
 FILLCELL_X32 FILLER_34_1 ();
 FILLCELL_X32 FILLER_34_33 ();
 FILLCELL_X32 FILLER_34_65 ();
 FILLCELL_X32 FILLER_34_97 ();
 FILLCELL_X32 FILLER_34_129 ();
 FILLCELL_X8 FILLER_34_161 ();
 FILLCELL_X2 FILLER_34_169 ();
 FILLCELL_X1 FILLER_34_171 ();
 FILLCELL_X4 FILLER_34_182 ();
 FILLCELL_X2 FILLER_34_186 ();
 FILLCELL_X1 FILLER_34_188 ();
 FILLCELL_X2 FILLER_34_217 ();
 FILLCELL_X2 FILLER_34_223 ();
 FILLCELL_X2 FILLER_34_229 ();
 FILLCELL_X2 FILLER_34_240 ();
 FILLCELL_X2 FILLER_34_259 ();
 FILLCELL_X4 FILLER_34_291 ();
 FILLCELL_X2 FILLER_34_295 ();
 FILLCELL_X1 FILLER_34_297 ();
 FILLCELL_X8 FILLER_34_301 ();
 FILLCELL_X2 FILLER_34_309 ();
 FILLCELL_X1 FILLER_34_311 ();
 FILLCELL_X2 FILLER_34_329 ();
 FILLCELL_X4 FILLER_34_338 ();
 FILLCELL_X2 FILLER_34_342 ();
 FILLCELL_X1 FILLER_34_361 ();
 FILLCELL_X16 FILLER_34_381 ();
 FILLCELL_X8 FILLER_34_397 ();
 FILLCELL_X4 FILLER_34_405 ();
 FILLCELL_X2 FILLER_34_409 ();
 FILLCELL_X1 FILLER_34_411 ();
 FILLCELL_X4 FILLER_34_429 ();
 FILLCELL_X2 FILLER_34_433 ();
 FILLCELL_X1 FILLER_34_435 ();
 FILLCELL_X4 FILLER_34_467 ();
 FILLCELL_X2 FILLER_34_471 ();
 FILLCELL_X1 FILLER_34_473 ();
 FILLCELL_X8 FILLER_34_484 ();
 FILLCELL_X4 FILLER_34_492 ();
 FILLCELL_X4 FILLER_34_513 ();
 FILLCELL_X1 FILLER_34_517 ();
 FILLCELL_X32 FILLER_34_542 ();
 FILLCELL_X8 FILLER_34_574 ();
 FILLCELL_X8 FILLER_34_591 ();
 FILLCELL_X1 FILLER_34_599 ();
 FILLCELL_X2 FILLER_34_629 ();
 FILLCELL_X2 FILLER_34_632 ();
 FILLCELL_X1 FILLER_34_634 ();
 FILLCELL_X8 FILLER_34_648 ();
 FILLCELL_X2 FILLER_34_656 ();
 FILLCELL_X16 FILLER_34_662 ();
 FILLCELL_X8 FILLER_34_678 ();
 FILLCELL_X2 FILLER_34_686 ();
 FILLCELL_X1 FILLER_34_688 ();
 FILLCELL_X32 FILLER_34_708 ();
 FILLCELL_X16 FILLER_34_740 ();
 FILLCELL_X2 FILLER_34_759 ();
 FILLCELL_X2 FILLER_34_776 ();
 FILLCELL_X1 FILLER_34_785 ();
 FILLCELL_X1 FILLER_34_817 ();
 FILLCELL_X2 FILLER_34_829 ();
 FILLCELL_X1 FILLER_34_831 ();
 FILLCELL_X4 FILLER_34_851 ();
 FILLCELL_X2 FILLER_34_855 ();
 FILLCELL_X1 FILLER_34_857 ();
 FILLCELL_X8 FILLER_34_862 ();
 FILLCELL_X8 FILLER_34_888 ();
 FILLCELL_X4 FILLER_34_896 ();
 FILLCELL_X4 FILLER_34_904 ();
 FILLCELL_X4 FILLER_34_927 ();
 FILLCELL_X1 FILLER_34_931 ();
 FILLCELL_X16 FILLER_34_939 ();
 FILLCELL_X2 FILLER_34_955 ();
 FILLCELL_X32 FILLER_34_976 ();
 FILLCELL_X8 FILLER_34_1008 ();
 FILLCELL_X4 FILLER_34_1033 ();
 FILLCELL_X2 FILLER_34_1037 ();
 FILLCELL_X2 FILLER_34_1084 ();
 FILLCELL_X8 FILLER_34_1107 ();
 FILLCELL_X1 FILLER_34_1115 ();
 FILLCELL_X1 FILLER_34_1138 ();
 FILLCELL_X2 FILLER_34_1166 ();
 FILLCELL_X4 FILLER_34_1175 ();
 FILLCELL_X4 FILLER_34_1187 ();
 FILLCELL_X8 FILLER_34_1198 ();
 FILLCELL_X2 FILLER_34_1206 ();
 FILLCELL_X1 FILLER_34_1208 ();
 FILLCELL_X32 FILLER_35_1 ();
 FILLCELL_X16 FILLER_35_33 ();
 FILLCELL_X4 FILLER_35_49 ();
 FILLCELL_X2 FILLER_35_53 ();
 FILLCELL_X32 FILLER_35_72 ();
 FILLCELL_X16 FILLER_35_104 ();
 FILLCELL_X8 FILLER_35_120 ();
 FILLCELL_X4 FILLER_35_128 ();
 FILLCELL_X32 FILLER_35_136 ();
 FILLCELL_X32 FILLER_35_168 ();
 FILLCELL_X2 FILLER_35_200 ();
 FILLCELL_X2 FILLER_35_212 ();
 FILLCELL_X1 FILLER_35_214 ();
 FILLCELL_X8 FILLER_35_232 ();
 FILLCELL_X4 FILLER_35_240 ();
 FILLCELL_X8 FILLER_35_274 ();
 FILLCELL_X2 FILLER_35_282 ();
 FILLCELL_X1 FILLER_35_284 ();
 FILLCELL_X8 FILLER_35_290 ();
 FILLCELL_X4 FILLER_35_315 ();
 FILLCELL_X2 FILLER_35_319 ();
 FILLCELL_X1 FILLER_35_321 ();
 FILLCELL_X1 FILLER_35_335 ();
 FILLCELL_X4 FILLER_35_389 ();
 FILLCELL_X2 FILLER_35_393 ();
 FILLCELL_X1 FILLER_35_420 ();
 FILLCELL_X4 FILLER_35_438 ();
 FILLCELL_X8 FILLER_35_447 ();
 FILLCELL_X4 FILLER_35_455 ();
 FILLCELL_X2 FILLER_35_459 ();
 FILLCELL_X1 FILLER_35_480 ();
 FILLCELL_X16 FILLER_35_500 ();
 FILLCELL_X2 FILLER_35_533 ();
 FILLCELL_X2 FILLER_35_544 ();
 FILLCELL_X1 FILLER_35_546 ();
 FILLCELL_X16 FILLER_35_556 ();
 FILLCELL_X16 FILLER_35_593 ();
 FILLCELL_X2 FILLER_35_609 ();
 FILLCELL_X2 FILLER_35_632 ();
 FILLCELL_X2 FILLER_35_647 ();
 FILLCELL_X1 FILLER_35_649 ();
 FILLCELL_X8 FILLER_35_659 ();
 FILLCELL_X1 FILLER_35_667 ();
 FILLCELL_X8 FILLER_35_678 ();
 FILLCELL_X4 FILLER_35_686 ();
 FILLCELL_X16 FILLER_35_699 ();
 FILLCELL_X4 FILLER_35_715 ();
 FILLCELL_X2 FILLER_35_719 ();
 FILLCELL_X1 FILLER_35_721 ();
 FILLCELL_X2 FILLER_35_739 ();
 FILLCELL_X1 FILLER_35_762 ();
 FILLCELL_X2 FILLER_35_768 ();
 FILLCELL_X2 FILLER_35_773 ();
 FILLCELL_X2 FILLER_35_790 ();
 FILLCELL_X1 FILLER_35_792 ();
 FILLCELL_X4 FILLER_35_857 ();
 FILLCELL_X8 FILLER_35_865 ();
 FILLCELL_X1 FILLER_35_873 ();
 FILLCELL_X2 FILLER_35_878 ();
 FILLCELL_X1 FILLER_35_880 ();
 FILLCELL_X1 FILLER_35_892 ();
 FILLCELL_X4 FILLER_35_921 ();
 FILLCELL_X2 FILLER_35_925 ();
 FILLCELL_X32 FILLER_35_931 ();
 FILLCELL_X32 FILLER_35_963 ();
 FILLCELL_X8 FILLER_35_995 ();
 FILLCELL_X4 FILLER_35_1003 ();
 FILLCELL_X2 FILLER_35_1007 ();
 FILLCELL_X1 FILLER_35_1023 ();
 FILLCELL_X4 FILLER_35_1031 ();
 FILLCELL_X2 FILLER_35_1035 ();
 FILLCELL_X2 FILLER_35_1057 ();
 FILLCELL_X4 FILLER_35_1097 ();
 FILLCELL_X8 FILLER_35_1108 ();
 FILLCELL_X1 FILLER_35_1116 ();
 FILLCELL_X2 FILLER_35_1122 ();
 FILLCELL_X1 FILLER_35_1124 ();
 FILLCELL_X4 FILLER_35_1133 ();
 FILLCELL_X1 FILLER_35_1137 ();
 FILLCELL_X1 FILLER_35_1154 ();
 FILLCELL_X1 FILLER_35_1160 ();
 FILLCELL_X2 FILLER_35_1171 ();
 FILLCELL_X1 FILLER_35_1184 ();
 FILLCELL_X2 FILLER_35_1190 ();
 FILLCELL_X4 FILLER_35_1202 ();
 FILLCELL_X2 FILLER_35_1206 ();
 FILLCELL_X1 FILLER_35_1208 ();
 FILLCELL_X32 FILLER_36_1 ();
 FILLCELL_X32 FILLER_36_33 ();
 FILLCELL_X16 FILLER_36_65 ();
 FILLCELL_X4 FILLER_36_81 ();
 FILLCELL_X2 FILLER_36_85 ();
 FILLCELL_X1 FILLER_36_100 ();
 FILLCELL_X8 FILLER_36_108 ();
 FILLCELL_X4 FILLER_36_156 ();
 FILLCELL_X4 FILLER_36_170 ();
 FILLCELL_X1 FILLER_36_174 ();
 FILLCELL_X8 FILLER_36_184 ();
 FILLCELL_X4 FILLER_36_192 ();
 FILLCELL_X2 FILLER_36_196 ();
 FILLCELL_X4 FILLER_36_210 ();
 FILLCELL_X1 FILLER_36_214 ();
 FILLCELL_X16 FILLER_36_222 ();
 FILLCELL_X2 FILLER_36_238 ();
 FILLCELL_X1 FILLER_36_240 ();
 FILLCELL_X2 FILLER_36_258 ();
 FILLCELL_X8 FILLER_36_265 ();
 FILLCELL_X32 FILLER_36_282 ();
 FILLCELL_X32 FILLER_36_314 ();
 FILLCELL_X4 FILLER_36_346 ();
 FILLCELL_X1 FILLER_36_350 ();
 FILLCELL_X4 FILLER_36_357 ();
 FILLCELL_X16 FILLER_36_363 ();
 FILLCELL_X16 FILLER_36_382 ();
 FILLCELL_X4 FILLER_36_398 ();
 FILLCELL_X2 FILLER_36_402 ();
 FILLCELL_X16 FILLER_36_411 ();
 FILLCELL_X16 FILLER_36_434 ();
 FILLCELL_X2 FILLER_36_450 ();
 FILLCELL_X4 FILLER_36_479 ();
 FILLCELL_X2 FILLER_36_483 ();
 FILLCELL_X16 FILLER_36_498 ();
 FILLCELL_X4 FILLER_36_514 ();
 FILLCELL_X2 FILLER_36_518 ();
 FILLCELL_X1 FILLER_36_520 ();
 FILLCELL_X1 FILLER_36_528 ();
 FILLCELL_X2 FILLER_36_543 ();
 FILLCELL_X1 FILLER_36_545 ();
 FILLCELL_X8 FILLER_36_550 ();
 FILLCELL_X2 FILLER_36_558 ();
 FILLCELL_X8 FILLER_36_601 ();
 FILLCELL_X4 FILLER_36_609 ();
 FILLCELL_X2 FILLER_36_613 ();
 FILLCELL_X1 FILLER_36_615 ();
 FILLCELL_X4 FILLER_36_625 ();
 FILLCELL_X2 FILLER_36_629 ();
 FILLCELL_X16 FILLER_36_645 ();
 FILLCELL_X8 FILLER_36_661 ();
 FILLCELL_X1 FILLER_36_669 ();
 FILLCELL_X16 FILLER_36_679 ();
 FILLCELL_X2 FILLER_36_712 ();
 FILLCELL_X1 FILLER_36_714 ();
 FILLCELL_X1 FILLER_36_744 ();
 FILLCELL_X1 FILLER_36_785 ();
 FILLCELL_X8 FILLER_36_836 ();
 FILLCELL_X4 FILLER_36_844 ();
 FILLCELL_X2 FILLER_36_848 ();
 FILLCELL_X1 FILLER_36_850 ();
 FILLCELL_X1 FILLER_36_869 ();
 FILLCELL_X4 FILLER_36_875 ();
 FILLCELL_X1 FILLER_36_879 ();
 FILLCELL_X2 FILLER_36_884 ();
 FILLCELL_X4 FILLER_36_905 ();
 FILLCELL_X2 FILLER_36_909 ();
 FILLCELL_X2 FILLER_36_915 ();
 FILLCELL_X1 FILLER_36_917 ();
 FILLCELL_X16 FILLER_36_938 ();
 FILLCELL_X8 FILLER_36_954 ();
 FILLCELL_X2 FILLER_36_962 ();
 FILLCELL_X16 FILLER_36_987 ();
 FILLCELL_X8 FILLER_36_1003 ();
 FILLCELL_X2 FILLER_36_1011 ();
 FILLCELL_X1 FILLER_36_1013 ();
 FILLCELL_X1 FILLER_36_1030 ();
 FILLCELL_X1 FILLER_36_1052 ();
 FILLCELL_X4 FILLER_36_1090 ();
 FILLCELL_X2 FILLER_36_1094 ();
 FILLCELL_X1 FILLER_36_1096 ();
 FILLCELL_X8 FILLER_36_1112 ();
 FILLCELL_X2 FILLER_36_1120 ();
 FILLCELL_X1 FILLER_36_1122 ();
 FILLCELL_X2 FILLER_36_1127 ();
 FILLCELL_X2 FILLER_36_1133 ();
 FILLCELL_X2 FILLER_36_1138 ();
 FILLCELL_X2 FILLER_36_1144 ();
 FILLCELL_X1 FILLER_36_1154 ();
 FILLCELL_X1 FILLER_36_1159 ();
 FILLCELL_X1 FILLER_36_1163 ();
 FILLCELL_X2 FILLER_36_1178 ();
 FILLCELL_X2 FILLER_36_1187 ();
 FILLCELL_X8 FILLER_36_1199 ();
 FILLCELL_X2 FILLER_36_1207 ();
 FILLCELL_X32 FILLER_37_1 ();
 FILLCELL_X32 FILLER_37_33 ();
 FILLCELL_X16 FILLER_37_65 ();
 FILLCELL_X8 FILLER_37_81 ();
 FILLCELL_X2 FILLER_37_89 ();
 FILLCELL_X2 FILLER_37_109 ();
 FILLCELL_X1 FILLER_37_111 ();
 FILLCELL_X1 FILLER_37_147 ();
 FILLCELL_X2 FILLER_37_173 ();
 FILLCELL_X1 FILLER_37_175 ();
 FILLCELL_X2 FILLER_37_180 ();
 FILLCELL_X8 FILLER_37_189 ();
 FILLCELL_X4 FILLER_37_197 ();
 FILLCELL_X2 FILLER_37_201 ();
 FILLCELL_X8 FILLER_37_207 ();
 FILLCELL_X16 FILLER_37_232 ();
 FILLCELL_X8 FILLER_37_248 ();
 FILLCELL_X2 FILLER_37_256 ();
 FILLCELL_X32 FILLER_37_275 ();
 FILLCELL_X8 FILLER_37_307 ();
 FILLCELL_X2 FILLER_37_325 ();
 FILLCELL_X2 FILLER_37_331 ();
 FILLCELL_X1 FILLER_37_333 ();
 FILLCELL_X16 FILLER_37_348 ();
 FILLCELL_X8 FILLER_37_364 ();
 FILLCELL_X8 FILLER_37_382 ();
 FILLCELL_X4 FILLER_37_390 ();
 FILLCELL_X2 FILLER_37_394 ();
 FILLCELL_X32 FILLER_37_403 ();
 FILLCELL_X16 FILLER_37_435 ();
 FILLCELL_X8 FILLER_37_451 ();
 FILLCELL_X4 FILLER_37_459 ();
 FILLCELL_X1 FILLER_37_463 ();
 FILLCELL_X4 FILLER_37_467 ();
 FILLCELL_X4 FILLER_37_477 ();
 FILLCELL_X2 FILLER_37_481 ();
 FILLCELL_X1 FILLER_37_483 ();
 FILLCELL_X32 FILLER_37_498 ();
 FILLCELL_X2 FILLER_37_530 ();
 FILLCELL_X1 FILLER_37_532 ();
 FILLCELL_X16 FILLER_37_551 ();
 FILLCELL_X1 FILLER_37_567 ();
 FILLCELL_X4 FILLER_37_603 ();
 FILLCELL_X2 FILLER_37_626 ();
 FILLCELL_X1 FILLER_37_628 ();
 FILLCELL_X8 FILLER_37_648 ();
 FILLCELL_X1 FILLER_37_656 ();
 FILLCELL_X4 FILLER_37_674 ();
 FILLCELL_X2 FILLER_37_678 ();
 FILLCELL_X4 FILLER_37_697 ();
 FILLCELL_X2 FILLER_37_701 ();
 FILLCELL_X2 FILLER_37_729 ();
 FILLCELL_X2 FILLER_37_748 ();
 FILLCELL_X1 FILLER_37_750 ();
 FILLCELL_X1 FILLER_37_772 ();
 FILLCELL_X1 FILLER_37_792 ();
 FILLCELL_X8 FILLER_37_835 ();
 FILLCELL_X1 FILLER_37_843 ();
 FILLCELL_X4 FILLER_37_848 ();
 FILLCELL_X4 FILLER_37_859 ();
 FILLCELL_X1 FILLER_37_863 ();
 FILLCELL_X4 FILLER_37_886 ();
 FILLCELL_X1 FILLER_37_890 ();
 FILLCELL_X4 FILLER_37_894 ();
 FILLCELL_X1 FILLER_37_898 ();
 FILLCELL_X2 FILLER_37_903 ();
 FILLCELL_X1 FILLER_37_905 ();
 FILLCELL_X2 FILLER_37_922 ();
 FILLCELL_X1 FILLER_37_924 ();
 FILLCELL_X1 FILLER_37_933 ();
 FILLCELL_X2 FILLER_37_939 ();
 FILLCELL_X4 FILLER_37_946 ();
 FILLCELL_X2 FILLER_37_967 ();
 FILLCELL_X1 FILLER_37_969 ();
 FILLCELL_X2 FILLER_37_977 ();
 FILLCELL_X1 FILLER_37_979 ();
 FILLCELL_X16 FILLER_37_984 ();
 FILLCELL_X8 FILLER_37_1000 ();
 FILLCELL_X4 FILLER_37_1008 ();
 FILLCELL_X1 FILLER_37_1012 ();
 FILLCELL_X4 FILLER_37_1042 ();
 FILLCELL_X1 FILLER_37_1059 ();
 FILLCELL_X2 FILLER_37_1070 ();
 FILLCELL_X4 FILLER_37_1080 ();
 FILLCELL_X2 FILLER_37_1084 ();
 FILLCELL_X2 FILLER_37_1103 ();
 FILLCELL_X1 FILLER_37_1105 ();
 FILLCELL_X2 FILLER_37_1114 ();
 FILLCELL_X1 FILLER_37_1116 ();
 FILLCELL_X2 FILLER_37_1120 ();
 FILLCELL_X1 FILLER_37_1122 ();
 FILLCELL_X4 FILLER_37_1131 ();
 FILLCELL_X2 FILLER_37_1135 ();
 FILLCELL_X1 FILLER_37_1144 ();
 FILLCELL_X2 FILLER_37_1150 ();
 FILLCELL_X1 FILLER_37_1152 ();
 FILLCELL_X2 FILLER_37_1169 ();
 FILLCELL_X2 FILLER_37_1190 ();
 FILLCELL_X8 FILLER_37_1199 ();
 FILLCELL_X2 FILLER_37_1207 ();
 FILLCELL_X32 FILLER_38_1 ();
 FILLCELL_X32 FILLER_38_33 ();
 FILLCELL_X1 FILLER_38_65 ();
 FILLCELL_X1 FILLER_38_97 ();
 FILLCELL_X2 FILLER_38_105 ();
 FILLCELL_X2 FILLER_38_114 ();
 FILLCELL_X2 FILLER_38_123 ();
 FILLCELL_X4 FILLER_38_158 ();
 FILLCELL_X2 FILLER_38_162 ();
 FILLCELL_X1 FILLER_38_164 ();
 FILLCELL_X8 FILLER_38_168 ();
 FILLCELL_X4 FILLER_38_176 ();
 FILLCELL_X1 FILLER_38_180 ();
 FILLCELL_X8 FILLER_38_186 ();
 FILLCELL_X1 FILLER_38_199 ();
 FILLCELL_X2 FILLER_38_210 ();
 FILLCELL_X1 FILLER_38_212 ();
 FILLCELL_X8 FILLER_38_222 ();
 FILLCELL_X2 FILLER_38_230 ();
 FILLCELL_X16 FILLER_38_237 ();
 FILLCELL_X8 FILLER_38_253 ();
 FILLCELL_X1 FILLER_38_261 ();
 FILLCELL_X4 FILLER_38_267 ();
 FILLCELL_X2 FILLER_38_271 ();
 FILLCELL_X1 FILLER_38_273 ();
 FILLCELL_X1 FILLER_38_323 ();
 FILLCELL_X8 FILLER_38_334 ();
 FILLCELL_X2 FILLER_38_342 ();
 FILLCELL_X4 FILLER_38_351 ();
 FILLCELL_X2 FILLER_38_355 ();
 FILLCELL_X2 FILLER_38_375 ();
 FILLCELL_X1 FILLER_38_377 ();
 FILLCELL_X4 FILLER_38_381 ();
 FILLCELL_X1 FILLER_38_385 ();
 FILLCELL_X4 FILLER_38_396 ();
 FILLCELL_X4 FILLER_38_421 ();
 FILLCELL_X2 FILLER_38_432 ();
 FILLCELL_X8 FILLER_38_447 ();
 FILLCELL_X4 FILLER_38_455 ();
 FILLCELL_X2 FILLER_38_459 ();
 FILLCELL_X1 FILLER_38_487 ();
 FILLCELL_X8 FILLER_38_494 ();
 FILLCELL_X4 FILLER_38_502 ();
 FILLCELL_X1 FILLER_38_506 ();
 FILLCELL_X4 FILLER_38_524 ();
 FILLCELL_X2 FILLER_38_528 ();
 FILLCELL_X8 FILLER_38_550 ();
 FILLCELL_X4 FILLER_38_558 ();
 FILLCELL_X2 FILLER_38_562 ();
 FILLCELL_X1 FILLER_38_564 ();
 FILLCELL_X2 FILLER_38_611 ();
 FILLCELL_X8 FILLER_38_651 ();
 FILLCELL_X4 FILLER_38_659 ();
 FILLCELL_X1 FILLER_38_663 ();
 FILLCELL_X16 FILLER_38_712 ();
 FILLCELL_X8 FILLER_38_728 ();
 FILLCELL_X2 FILLER_38_736 ();
 FILLCELL_X1 FILLER_38_738 ();
 FILLCELL_X4 FILLER_38_762 ();
 FILLCELL_X1 FILLER_38_766 ();
 FILLCELL_X2 FILLER_38_786 ();
 FILLCELL_X2 FILLER_38_802 ();
 FILLCELL_X1 FILLER_38_859 ();
 FILLCELL_X1 FILLER_38_878 ();
 FILLCELL_X4 FILLER_38_914 ();
 FILLCELL_X1 FILLER_38_918 ();
 FILLCELL_X4 FILLER_38_925 ();
 FILLCELL_X2 FILLER_38_934 ();
 FILLCELL_X32 FILLER_38_945 ();
 FILLCELL_X32 FILLER_38_977 ();
 FILLCELL_X4 FILLER_38_1009 ();
 FILLCELL_X8 FILLER_38_1023 ();
 FILLCELL_X4 FILLER_38_1031 ();
 FILLCELL_X4 FILLER_38_1053 ();
 FILLCELL_X8 FILLER_38_1060 ();
 FILLCELL_X1 FILLER_38_1068 ();
 FILLCELL_X4 FILLER_38_1081 ();
 FILLCELL_X4 FILLER_38_1089 ();
 FILLCELL_X4 FILLER_38_1097 ();
 FILLCELL_X2 FILLER_38_1122 ();
 FILLCELL_X1 FILLER_38_1124 ();
 FILLCELL_X1 FILLER_38_1128 ();
 FILLCELL_X4 FILLER_38_1140 ();
 FILLCELL_X1 FILLER_38_1144 ();
 FILLCELL_X4 FILLER_38_1149 ();
 FILLCELL_X2 FILLER_38_1153 ();
 FILLCELL_X1 FILLER_38_1155 ();
 FILLCELL_X4 FILLER_38_1183 ();
 FILLCELL_X2 FILLER_38_1187 ();
 FILLCELL_X16 FILLER_38_1192 ();
 FILLCELL_X1 FILLER_38_1208 ();
 FILLCELL_X32 FILLER_39_1 ();
 FILLCELL_X32 FILLER_39_33 ();
 FILLCELL_X4 FILLER_39_65 ();
 FILLCELL_X2 FILLER_39_69 ();
 FILLCELL_X1 FILLER_39_71 ();
 FILLCELL_X2 FILLER_39_110 ();
 FILLCELL_X2 FILLER_39_123 ();
 FILLCELL_X1 FILLER_39_125 ();
 FILLCELL_X1 FILLER_39_141 ();
 FILLCELL_X2 FILLER_39_159 ();
 FILLCELL_X1 FILLER_39_169 ();
 FILLCELL_X8 FILLER_39_178 ();
 FILLCELL_X1 FILLER_39_186 ();
 FILLCELL_X1 FILLER_39_194 ();
 FILLCELL_X4 FILLER_39_202 ();
 FILLCELL_X1 FILLER_39_206 ();
 FILLCELL_X32 FILLER_39_225 ();
 FILLCELL_X16 FILLER_39_257 ();
 FILLCELL_X2 FILLER_39_273 ();
 FILLCELL_X1 FILLER_39_275 ();
 FILLCELL_X2 FILLER_39_296 ();
 FILLCELL_X1 FILLER_39_309 ();
 FILLCELL_X8 FILLER_39_341 ();
 FILLCELL_X4 FILLER_39_349 ();
 FILLCELL_X2 FILLER_39_353 ();
 FILLCELL_X1 FILLER_39_372 ();
 FILLCELL_X4 FILLER_39_390 ();
 FILLCELL_X16 FILLER_39_437 ();
 FILLCELL_X2 FILLER_39_453 ();
 FILLCELL_X4 FILLER_39_460 ();
 FILLCELL_X2 FILLER_39_494 ();
 FILLCELL_X1 FILLER_39_496 ();
 FILLCELL_X2 FILLER_39_503 ();
 FILLCELL_X1 FILLER_39_505 ();
 FILLCELL_X4 FILLER_39_526 ();
 FILLCELL_X1 FILLER_39_530 ();
 FILLCELL_X4 FILLER_39_536 ();
 FILLCELL_X1 FILLER_39_550 ();
 FILLCELL_X4 FILLER_39_557 ();
 FILLCELL_X2 FILLER_39_561 ();
 FILLCELL_X1 FILLER_39_566 ();
 FILLCELL_X2 FILLER_39_574 ();
 FILLCELL_X2 FILLER_39_582 ();
 FILLCELL_X8 FILLER_39_590 ();
 FILLCELL_X4 FILLER_39_607 ();
 FILLCELL_X8 FILLER_39_615 ();
 FILLCELL_X4 FILLER_39_623 ();
 FILLCELL_X2 FILLER_39_627 ();
 FILLCELL_X4 FILLER_39_653 ();
 FILLCELL_X4 FILLER_39_674 ();
 FILLCELL_X2 FILLER_39_678 ();
 FILLCELL_X1 FILLER_39_688 ();
 FILLCELL_X1 FILLER_39_696 ();
 FILLCELL_X1 FILLER_39_704 ();
 FILLCELL_X16 FILLER_39_711 ();
 FILLCELL_X8 FILLER_39_727 ();
 FILLCELL_X4 FILLER_39_735 ();
 FILLCELL_X2 FILLER_39_739 ();
 FILLCELL_X1 FILLER_39_741 ();
 FILLCELL_X4 FILLER_39_763 ();
 FILLCELL_X1 FILLER_39_767 ();
 FILLCELL_X2 FILLER_39_781 ();
 FILLCELL_X1 FILLER_39_794 ();
 FILLCELL_X4 FILLER_39_835 ();
 FILLCELL_X2 FILLER_39_839 ();
 FILLCELL_X1 FILLER_39_841 ();
 FILLCELL_X16 FILLER_39_857 ();
 FILLCELL_X8 FILLER_39_873 ();
 FILLCELL_X4 FILLER_39_881 ();
 FILLCELL_X8 FILLER_39_888 ();
 FILLCELL_X4 FILLER_39_896 ();
 FILLCELL_X4 FILLER_39_904 ();
 FILLCELL_X1 FILLER_39_908 ();
 FILLCELL_X2 FILLER_39_913 ();
 FILLCELL_X32 FILLER_39_925 ();
 FILLCELL_X32 FILLER_39_957 ();
 FILLCELL_X16 FILLER_39_989 ();
 FILLCELL_X8 FILLER_39_1005 ();
 FILLCELL_X4 FILLER_39_1013 ();
 FILLCELL_X2 FILLER_39_1017 ();
 FILLCELL_X1 FILLER_39_1019 ();
 FILLCELL_X1 FILLER_39_1027 ();
 FILLCELL_X2 FILLER_39_1032 ();
 FILLCELL_X2 FILLER_39_1064 ();
 FILLCELL_X4 FILLER_39_1089 ();
 FILLCELL_X4 FILLER_39_1097 ();
 FILLCELL_X1 FILLER_39_1101 ();
 FILLCELL_X2 FILLER_39_1118 ();
 FILLCELL_X1 FILLER_39_1120 ();
 FILLCELL_X2 FILLER_39_1125 ();
 FILLCELL_X2 FILLER_39_1140 ();
 FILLCELL_X4 FILLER_39_1160 ();
 FILLCELL_X4 FILLER_39_1168 ();
 FILLCELL_X2 FILLER_39_1176 ();
 FILLCELL_X1 FILLER_39_1178 ();
 FILLCELL_X16 FILLER_39_1184 ();
 FILLCELL_X8 FILLER_39_1200 ();
 FILLCELL_X1 FILLER_39_1208 ();
 FILLCELL_X32 FILLER_40_1 ();
 FILLCELL_X16 FILLER_40_33 ();
 FILLCELL_X8 FILLER_40_49 ();
 FILLCELL_X4 FILLER_40_57 ();
 FILLCELL_X2 FILLER_40_61 ();
 FILLCELL_X2 FILLER_40_92 ();
 FILLCELL_X1 FILLER_40_131 ();
 FILLCELL_X2 FILLER_40_136 ();
 FILLCELL_X1 FILLER_40_138 ();
 FILLCELL_X2 FILLER_40_143 ();
 FILLCELL_X1 FILLER_40_152 ();
 FILLCELL_X2 FILLER_40_157 ();
 FILLCELL_X4 FILLER_40_173 ();
 FILLCELL_X2 FILLER_40_177 ();
 FILLCELL_X1 FILLER_40_179 ();
 FILLCELL_X1 FILLER_40_189 ();
 FILLCELL_X32 FILLER_40_230 ();
 FILLCELL_X1 FILLER_40_285 ();
 FILLCELL_X1 FILLER_40_307 ();
 FILLCELL_X2 FILLER_40_341 ();
 FILLCELL_X1 FILLER_40_343 ();
 FILLCELL_X4 FILLER_40_351 ();
 FILLCELL_X2 FILLER_40_370 ();
 FILLCELL_X1 FILLER_40_372 ();
 FILLCELL_X1 FILLER_40_377 ();
 FILLCELL_X4 FILLER_40_388 ();
 FILLCELL_X2 FILLER_40_392 ();
 FILLCELL_X1 FILLER_40_394 ();
 FILLCELL_X4 FILLER_40_406 ();
 FILLCELL_X1 FILLER_40_435 ();
 FILLCELL_X4 FILLER_40_455 ();
 FILLCELL_X2 FILLER_40_459 ();
 FILLCELL_X1 FILLER_40_483 ();
 FILLCELL_X4 FILLER_40_530 ();
 FILLCELL_X2 FILLER_40_551 ();
 FILLCELL_X1 FILLER_40_553 ();
 FILLCELL_X2 FILLER_40_573 ();
 FILLCELL_X1 FILLER_40_575 ();
 FILLCELL_X2 FILLER_40_582 ();
 FILLCELL_X1 FILLER_40_584 ();
 FILLCELL_X2 FILLER_40_594 ();
 FILLCELL_X1 FILLER_40_596 ();
 FILLCELL_X4 FILLER_40_607 ();
 FILLCELL_X1 FILLER_40_611 ();
 FILLCELL_X8 FILLER_40_619 ();
 FILLCELL_X4 FILLER_40_627 ();
 FILLCELL_X1 FILLER_40_632 ();
 FILLCELL_X8 FILLER_40_655 ();
 FILLCELL_X4 FILLER_40_663 ();
 FILLCELL_X2 FILLER_40_676 ();
 FILLCELL_X1 FILLER_40_678 ();
 FILLCELL_X2 FILLER_40_685 ();
 FILLCELL_X1 FILLER_40_693 ();
 FILLCELL_X1 FILLER_40_698 ();
 FILLCELL_X8 FILLER_40_703 ();
 FILLCELL_X4 FILLER_40_711 ();
 FILLCELL_X8 FILLER_40_724 ();
 FILLCELL_X4 FILLER_40_732 ();
 FILLCELL_X2 FILLER_40_736 ();
 FILLCELL_X1 FILLER_40_738 ();
 FILLCELL_X2 FILLER_40_753 ();
 FILLCELL_X1 FILLER_40_755 ();
 FILLCELL_X2 FILLER_40_796 ();
 FILLCELL_X1 FILLER_40_848 ();
 FILLCELL_X2 FILLER_40_860 ();
 FILLCELL_X1 FILLER_40_865 ();
 FILLCELL_X2 FILLER_40_894 ();
 FILLCELL_X32 FILLER_40_934 ();
 FILLCELL_X4 FILLER_40_966 ();
 FILLCELL_X2 FILLER_40_970 ();
 FILLCELL_X8 FILLER_40_977 ();
 FILLCELL_X2 FILLER_40_985 ();
 FILLCELL_X1 FILLER_40_987 ();
 FILLCELL_X8 FILLER_40_1005 ();
 FILLCELL_X2 FILLER_40_1013 ();
 FILLCELL_X8 FILLER_40_1024 ();
 FILLCELL_X2 FILLER_40_1054 ();
 FILLCELL_X1 FILLER_40_1060 ();
 FILLCELL_X2 FILLER_40_1070 ();
 FILLCELL_X1 FILLER_40_1072 ();
 FILLCELL_X8 FILLER_40_1076 ();
 FILLCELL_X2 FILLER_40_1084 ();
 FILLCELL_X1 FILLER_40_1086 ();
 FILLCELL_X4 FILLER_40_1094 ();
 FILLCELL_X2 FILLER_40_1098 ();
 FILLCELL_X1 FILLER_40_1100 ();
 FILLCELL_X1 FILLER_40_1110 ();
 FILLCELL_X4 FILLER_40_1115 ();
 FILLCELL_X2 FILLER_40_1119 ();
 FILLCELL_X2 FILLER_40_1145 ();
 FILLCELL_X1 FILLER_40_1147 ();
 FILLCELL_X2 FILLER_40_1154 ();
 FILLCELL_X2 FILLER_40_1160 ();
 FILLCELL_X4 FILLER_40_1173 ();
 FILLCELL_X2 FILLER_40_1177 ();
 FILLCELL_X16 FILLER_40_1182 ();
 FILLCELL_X8 FILLER_40_1198 ();
 FILLCELL_X2 FILLER_40_1206 ();
 FILLCELL_X1 FILLER_40_1208 ();
 FILLCELL_X32 FILLER_41_1 ();
 FILLCELL_X16 FILLER_41_33 ();
 FILLCELL_X4 FILLER_41_49 ();
 FILLCELL_X2 FILLER_41_103 ();
 FILLCELL_X2 FILLER_41_112 ();
 FILLCELL_X1 FILLER_41_122 ();
 FILLCELL_X2 FILLER_41_127 ();
 FILLCELL_X1 FILLER_41_129 ();
 FILLCELL_X1 FILLER_41_145 ();
 FILLCELL_X2 FILLER_41_153 ();
 FILLCELL_X1 FILLER_41_155 ();
 FILLCELL_X4 FILLER_41_165 ();
 FILLCELL_X1 FILLER_41_177 ();
 FILLCELL_X1 FILLER_41_182 ();
 FILLCELL_X2 FILLER_41_195 ();
 FILLCELL_X1 FILLER_41_197 ();
 FILLCELL_X2 FILLER_41_205 ();
 FILLCELL_X4 FILLER_41_236 ();
 FILLCELL_X2 FILLER_41_240 ();
 FILLCELL_X8 FILLER_41_255 ();
 FILLCELL_X4 FILLER_41_263 ();
 FILLCELL_X1 FILLER_41_267 ();
 FILLCELL_X1 FILLER_41_313 ();
 FILLCELL_X4 FILLER_41_325 ();
 FILLCELL_X2 FILLER_41_329 ();
 FILLCELL_X1 FILLER_41_335 ();
 FILLCELL_X8 FILLER_41_340 ();
 FILLCELL_X2 FILLER_41_348 ();
 FILLCELL_X4 FILLER_41_361 ();
 FILLCELL_X4 FILLER_41_387 ();
 FILLCELL_X2 FILLER_41_405 ();
 FILLCELL_X4 FILLER_41_411 ();
 FILLCELL_X1 FILLER_41_415 ();
 FILLCELL_X32 FILLER_41_424 ();
 FILLCELL_X4 FILLER_41_456 ();
 FILLCELL_X1 FILLER_41_460 ();
 FILLCELL_X1 FILLER_41_474 ();
 FILLCELL_X1 FILLER_41_485 ();
 FILLCELL_X8 FILLER_41_510 ();
 FILLCELL_X4 FILLER_41_518 ();
 FILLCELL_X2 FILLER_41_522 ();
 FILLCELL_X1 FILLER_41_524 ();
 FILLCELL_X4 FILLER_41_542 ();
 FILLCELL_X2 FILLER_41_546 ();
 FILLCELL_X1 FILLER_41_555 ();
 FILLCELL_X8 FILLER_41_566 ();
 FILLCELL_X1 FILLER_41_574 ();
 FILLCELL_X2 FILLER_41_596 ();
 FILLCELL_X16 FILLER_41_604 ();
 FILLCELL_X8 FILLER_41_620 ();
 FILLCELL_X1 FILLER_41_628 ();
 FILLCELL_X1 FILLER_41_635 ();
 FILLCELL_X2 FILLER_41_645 ();
 FILLCELL_X1 FILLER_41_647 ();
 FILLCELL_X1 FILLER_41_670 ();
 FILLCELL_X4 FILLER_41_685 ();
 FILLCELL_X1 FILLER_41_695 ();
 FILLCELL_X2 FILLER_41_702 ();
 FILLCELL_X1 FILLER_41_704 ();
 FILLCELL_X32 FILLER_41_724 ();
 FILLCELL_X1 FILLER_41_786 ();
 FILLCELL_X8 FILLER_41_815 ();
 FILLCELL_X4 FILLER_41_823 ();
 FILLCELL_X2 FILLER_41_827 ();
 FILLCELL_X1 FILLER_41_840 ();
 FILLCELL_X2 FILLER_41_869 ();
 FILLCELL_X1 FILLER_41_917 ();
 FILLCELL_X16 FILLER_41_928 ();
 FILLCELL_X4 FILLER_41_944 ();
 FILLCELL_X2 FILLER_41_948 ();
 FILLCELL_X16 FILLER_41_967 ();
 FILLCELL_X4 FILLER_41_992 ();
 FILLCELL_X2 FILLER_41_996 ();
 FILLCELL_X1 FILLER_41_1055 ();
 FILLCELL_X2 FILLER_41_1068 ();
 FILLCELL_X8 FILLER_41_1074 ();
 FILLCELL_X2 FILLER_41_1082 ();
 FILLCELL_X1 FILLER_41_1084 ();
 FILLCELL_X1 FILLER_41_1105 ();
 FILLCELL_X2 FILLER_41_1117 ();
 FILLCELL_X1 FILLER_41_1123 ();
 FILLCELL_X1 FILLER_41_1127 ();
 FILLCELL_X2 FILLER_41_1157 ();
 FILLCELL_X1 FILLER_41_1159 ();
 FILLCELL_X2 FILLER_41_1168 ();
 FILLCELL_X1 FILLER_41_1174 ();
 FILLCELL_X16 FILLER_41_1192 ();
 FILLCELL_X1 FILLER_41_1208 ();
 FILLCELL_X8 FILLER_42_1 ();
 FILLCELL_X4 FILLER_42_9 ();
 FILLCELL_X1 FILLER_42_13 ();
 FILLCELL_X16 FILLER_42_31 ();
 FILLCELL_X2 FILLER_42_47 ();
 FILLCELL_X2 FILLER_42_70 ();
 FILLCELL_X2 FILLER_42_95 ();
 FILLCELL_X4 FILLER_42_119 ();
 FILLCELL_X2 FILLER_42_123 ();
 FILLCELL_X1 FILLER_42_125 ();
 FILLCELL_X1 FILLER_42_147 ();
 FILLCELL_X4 FILLER_42_159 ();
 FILLCELL_X1 FILLER_42_163 ();
 FILLCELL_X1 FILLER_42_167 ();
 FILLCELL_X2 FILLER_42_188 ();
 FILLCELL_X1 FILLER_42_190 ();
 FILLCELL_X2 FILLER_42_196 ();
 FILLCELL_X1 FILLER_42_213 ();
 FILLCELL_X16 FILLER_42_234 ();
 FILLCELL_X8 FILLER_42_250 ();
 FILLCELL_X2 FILLER_42_258 ();
 FILLCELL_X1 FILLER_42_260 ();
 FILLCELL_X8 FILLER_42_270 ();
 FILLCELL_X1 FILLER_42_278 ();
 FILLCELL_X4 FILLER_42_300 ();
 FILLCELL_X2 FILLER_42_304 ();
 FILLCELL_X1 FILLER_42_310 ();
 FILLCELL_X2 FILLER_42_323 ();
 FILLCELL_X1 FILLER_42_325 ();
 FILLCELL_X1 FILLER_42_341 ();
 FILLCELL_X1 FILLER_42_347 ();
 FILLCELL_X4 FILLER_42_351 ();
 FILLCELL_X2 FILLER_42_361 ();
 FILLCELL_X8 FILLER_42_371 ();
 FILLCELL_X1 FILLER_42_379 ();
 FILLCELL_X8 FILLER_42_384 ();
 FILLCELL_X4 FILLER_42_392 ();
 FILLCELL_X1 FILLER_42_396 ();
 FILLCELL_X4 FILLER_42_411 ();
 FILLCELL_X1 FILLER_42_415 ();
 FILLCELL_X4 FILLER_42_421 ();
 FILLCELL_X1 FILLER_42_425 ();
 FILLCELL_X16 FILLER_42_433 ();
 FILLCELL_X2 FILLER_42_449 ();
 FILLCELL_X1 FILLER_42_451 ();
 FILLCELL_X2 FILLER_42_469 ();
 FILLCELL_X4 FILLER_42_484 ();
 FILLCELL_X2 FILLER_42_488 ();
 FILLCELL_X4 FILLER_42_496 ();
 FILLCELL_X1 FILLER_42_500 ();
 FILLCELL_X4 FILLER_42_529 ();
 FILLCELL_X8 FILLER_42_542 ();
 FILLCELL_X1 FILLER_42_556 ();
 FILLCELL_X2 FILLER_42_559 ();
 FILLCELL_X1 FILLER_42_561 ();
 FILLCELL_X1 FILLER_42_565 ();
 FILLCELL_X8 FILLER_42_585 ();
 FILLCELL_X4 FILLER_42_593 ();
 FILLCELL_X1 FILLER_42_597 ();
 FILLCELL_X8 FILLER_42_620 ();
 FILLCELL_X2 FILLER_42_628 ();
 FILLCELL_X1 FILLER_42_630 ();
 FILLCELL_X8 FILLER_42_641 ();
 FILLCELL_X1 FILLER_42_649 ();
 FILLCELL_X1 FILLER_42_672 ();
 FILLCELL_X2 FILLER_42_679 ();
 FILLCELL_X1 FILLER_42_687 ();
 FILLCELL_X2 FILLER_42_694 ();
 FILLCELL_X8 FILLER_42_706 ();
 FILLCELL_X1 FILLER_42_714 ();
 FILLCELL_X16 FILLER_42_724 ();
 FILLCELL_X4 FILLER_42_740 ();
 FILLCELL_X1 FILLER_42_744 ();
 FILLCELL_X2 FILLER_42_754 ();
 FILLCELL_X4 FILLER_42_808 ();
 FILLCELL_X4 FILLER_42_816 ();
 FILLCELL_X2 FILLER_42_820 ();
 FILLCELL_X1 FILLER_42_822 ();
 FILLCELL_X4 FILLER_42_827 ();
 FILLCELL_X1 FILLER_42_831 ();
 FILLCELL_X4 FILLER_42_848 ();
 FILLCELL_X2 FILLER_42_852 ();
 FILLCELL_X2 FILLER_42_861 ();
 FILLCELL_X2 FILLER_42_883 ();
 FILLCELL_X8 FILLER_42_923 ();
 FILLCELL_X16 FILLER_42_942 ();
 FILLCELL_X4 FILLER_42_958 ();
 FILLCELL_X1 FILLER_42_962 ();
 FILLCELL_X8 FILLER_42_972 ();
 FILLCELL_X2 FILLER_42_980 ();
 FILLCELL_X8 FILLER_42_992 ();
 FILLCELL_X2 FILLER_42_1000 ();
 FILLCELL_X1 FILLER_42_1002 ();
 FILLCELL_X4 FILLER_42_1021 ();
 FILLCELL_X1 FILLER_42_1025 ();
 FILLCELL_X4 FILLER_42_1031 ();
 FILLCELL_X2 FILLER_42_1035 ();
 FILLCELL_X1 FILLER_42_1037 ();
 FILLCELL_X2 FILLER_42_1052 ();
 FILLCELL_X1 FILLER_42_1064 ();
 FILLCELL_X2 FILLER_42_1111 ();
 FILLCELL_X1 FILLER_42_1120 ();
 FILLCELL_X4 FILLER_42_1129 ();
 FILLCELL_X1 FILLER_42_1141 ();
 FILLCELL_X1 FILLER_42_1146 ();
 FILLCELL_X1 FILLER_42_1151 ();
 FILLCELL_X4 FILLER_42_1161 ();
 FILLCELL_X2 FILLER_42_1165 ();
 FILLCELL_X2 FILLER_42_1170 ();
 FILLCELL_X1 FILLER_42_1172 ();
 FILLCELL_X16 FILLER_42_1188 ();
 FILLCELL_X4 FILLER_42_1204 ();
 FILLCELL_X1 FILLER_42_1208 ();
 FILLCELL_X32 FILLER_43_1 ();
 FILLCELL_X16 FILLER_43_33 ();
 FILLCELL_X2 FILLER_43_49 ();
 FILLCELL_X1 FILLER_43_51 ();
 FILLCELL_X4 FILLER_43_104 ();
 FILLCELL_X2 FILLER_43_119 ();
 FILLCELL_X2 FILLER_43_136 ();
 FILLCELL_X1 FILLER_43_138 ();
 FILLCELL_X2 FILLER_43_154 ();
 FILLCELL_X8 FILLER_43_161 ();
 FILLCELL_X4 FILLER_43_169 ();
 FILLCELL_X2 FILLER_43_173 ();
 FILLCELL_X1 FILLER_43_179 ();
 FILLCELL_X2 FILLER_43_191 ();
 FILLCELL_X2 FILLER_43_202 ();
 FILLCELL_X1 FILLER_43_204 ();
 FILLCELL_X1 FILLER_43_208 ();
 FILLCELL_X1 FILLER_43_213 ();
 FILLCELL_X2 FILLER_43_218 ();
 FILLCELL_X1 FILLER_43_220 ();
 FILLCELL_X16 FILLER_43_238 ();
 FILLCELL_X8 FILLER_43_254 ();
 FILLCELL_X2 FILLER_43_262 ();
 FILLCELL_X1 FILLER_43_264 ();
 FILLCELL_X1 FILLER_43_293 ();
 FILLCELL_X2 FILLER_43_303 ();
 FILLCELL_X4 FILLER_43_322 ();
 FILLCELL_X2 FILLER_43_326 ();
 FILLCELL_X1 FILLER_43_328 ();
 FILLCELL_X2 FILLER_43_340 ();
 FILLCELL_X1 FILLER_43_342 ();
 FILLCELL_X2 FILLER_43_355 ();
 FILLCELL_X1 FILLER_43_357 ();
 FILLCELL_X1 FILLER_43_379 ();
 FILLCELL_X2 FILLER_43_389 ();
 FILLCELL_X2 FILLER_43_399 ();
 FILLCELL_X1 FILLER_43_405 ();
 FILLCELL_X1 FILLER_43_419 ();
 FILLCELL_X32 FILLER_43_431 ();
 FILLCELL_X2 FILLER_43_463 ();
 FILLCELL_X1 FILLER_43_477 ();
 FILLCELL_X16 FILLER_43_494 ();
 FILLCELL_X2 FILLER_43_510 ();
 FILLCELL_X8 FILLER_43_521 ();
 FILLCELL_X1 FILLER_43_529 ();
 FILLCELL_X4 FILLER_43_548 ();
 FILLCELL_X2 FILLER_43_552 ();
 FILLCELL_X1 FILLER_43_554 ();
 FILLCELL_X8 FILLER_43_570 ();
 FILLCELL_X4 FILLER_43_578 ();
 FILLCELL_X1 FILLER_43_582 ();
 FILLCELL_X1 FILLER_43_590 ();
 FILLCELL_X2 FILLER_43_601 ();
 FILLCELL_X1 FILLER_43_603 ();
 FILLCELL_X2 FILLER_43_618 ();
 FILLCELL_X4 FILLER_43_666 ();
 FILLCELL_X1 FILLER_43_670 ();
 FILLCELL_X2 FILLER_43_681 ();
 FILLCELL_X1 FILLER_43_683 ();
 FILLCELL_X2 FILLER_43_694 ();
 FILLCELL_X1 FILLER_43_696 ();
 FILLCELL_X2 FILLER_43_703 ();
 FILLCELL_X1 FILLER_43_705 ();
 FILLCELL_X32 FILLER_43_727 ();
 FILLCELL_X8 FILLER_43_769 ();
 FILLCELL_X1 FILLER_43_777 ();
 FILLCELL_X2 FILLER_43_798 ();
 FILLCELL_X1 FILLER_43_800 ();
 FILLCELL_X8 FILLER_43_827 ();
 FILLCELL_X1 FILLER_43_835 ();
 FILLCELL_X2 FILLER_43_854 ();
 FILLCELL_X2 FILLER_43_861 ();
 FILLCELL_X1 FILLER_43_863 ();
 FILLCELL_X2 FILLER_43_867 ();
 FILLCELL_X1 FILLER_43_869 ();
 FILLCELL_X2 FILLER_43_873 ();
 FILLCELL_X1 FILLER_43_875 ();
 FILLCELL_X8 FILLER_43_888 ();
 FILLCELL_X2 FILLER_43_907 ();
 FILLCELL_X4 FILLER_43_914 ();
 FILLCELL_X16 FILLER_43_951 ();
 FILLCELL_X4 FILLER_43_991 ();
 FILLCELL_X1 FILLER_43_995 ();
 FILLCELL_X8 FILLER_43_1009 ();
 FILLCELL_X1 FILLER_43_1017 ();
 FILLCELL_X2 FILLER_43_1022 ();
 FILLCELL_X8 FILLER_43_1044 ();
 FILLCELL_X4 FILLER_43_1052 ();
 FILLCELL_X2 FILLER_43_1060 ();
 FILLCELL_X1 FILLER_43_1062 ();
 FILLCELL_X1 FILLER_43_1072 ();
 FILLCELL_X1 FILLER_43_1088 ();
 FILLCELL_X8 FILLER_43_1109 ();
 FILLCELL_X1 FILLER_43_1117 ();
 FILLCELL_X8 FILLER_43_1121 ();
 FILLCELL_X1 FILLER_43_1129 ();
 FILLCELL_X4 FILLER_43_1143 ();
 FILLCELL_X2 FILLER_43_1149 ();
 FILLCELL_X4 FILLER_43_1170 ();
 FILLCELL_X2 FILLER_43_1184 ();
 FILLCELL_X1 FILLER_43_1186 ();
 FILLCELL_X16 FILLER_43_1191 ();
 FILLCELL_X2 FILLER_43_1207 ();
 FILLCELL_X32 FILLER_44_1 ();
 FILLCELL_X16 FILLER_44_33 ();
 FILLCELL_X8 FILLER_44_49 ();
 FILLCELL_X1 FILLER_44_57 ();
 FILLCELL_X2 FILLER_44_71 ();
 FILLCELL_X2 FILLER_44_84 ();
 FILLCELL_X16 FILLER_44_97 ();
 FILLCELL_X1 FILLER_44_113 ();
 FILLCELL_X4 FILLER_44_118 ();
 FILLCELL_X1 FILLER_44_122 ();
 FILLCELL_X1 FILLER_44_144 ();
 FILLCELL_X2 FILLER_44_149 ();
 FILLCELL_X1 FILLER_44_151 ();
 FILLCELL_X4 FILLER_44_203 ();
 FILLCELL_X2 FILLER_44_207 ();
 FILLCELL_X2 FILLER_44_213 ();
 FILLCELL_X32 FILLER_44_219 ();
 FILLCELL_X2 FILLER_44_251 ();
 FILLCELL_X1 FILLER_44_253 ();
 FILLCELL_X2 FILLER_44_284 ();
 FILLCELL_X1 FILLER_44_305 ();
 FILLCELL_X2 FILLER_44_313 ();
 FILLCELL_X2 FILLER_44_326 ();
 FILLCELL_X16 FILLER_44_341 ();
 FILLCELL_X4 FILLER_44_357 ();
 FILLCELL_X2 FILLER_44_383 ();
 FILLCELL_X1 FILLER_44_401 ();
 FILLCELL_X1 FILLER_44_407 ();
 FILLCELL_X2 FILLER_44_421 ();
 FILLCELL_X1 FILLER_44_423 ();
 FILLCELL_X16 FILLER_44_440 ();
 FILLCELL_X4 FILLER_44_456 ();
 FILLCELL_X2 FILLER_44_460 ();
 FILLCELL_X1 FILLER_44_462 ();
 FILLCELL_X4 FILLER_44_480 ();
 FILLCELL_X1 FILLER_44_547 ();
 FILLCELL_X4 FILLER_44_611 ();
 FILLCELL_X1 FILLER_44_630 ();
 FILLCELL_X2 FILLER_44_632 ();
 FILLCELL_X1 FILLER_44_634 ();
 FILLCELL_X16 FILLER_44_645 ();
 FILLCELL_X4 FILLER_44_661 ();
 FILLCELL_X16 FILLER_44_681 ();
 FILLCELL_X4 FILLER_44_706 ();
 FILLCELL_X2 FILLER_44_710 ();
 FILLCELL_X2 FILLER_44_718 ();
 FILLCELL_X1 FILLER_44_720 ();
 FILLCELL_X8 FILLER_44_741 ();
 FILLCELL_X2 FILLER_44_749 ();
 FILLCELL_X1 FILLER_44_751 ();
 FILLCELL_X2 FILLER_44_781 ();
 FILLCELL_X1 FILLER_44_800 ();
 FILLCELL_X2 FILLER_44_827 ();
 FILLCELL_X1 FILLER_44_864 ();
 FILLCELL_X8 FILLER_44_878 ();
 FILLCELL_X2 FILLER_44_886 ();
 FILLCELL_X1 FILLER_44_888 ();
 FILLCELL_X2 FILLER_44_898 ();
 FILLCELL_X4 FILLER_44_917 ();
 FILLCELL_X32 FILLER_44_932 ();
 FILLCELL_X16 FILLER_44_964 ();
 FILLCELL_X8 FILLER_44_980 ();
 FILLCELL_X2 FILLER_44_988 ();
 FILLCELL_X1 FILLER_44_990 ();
 FILLCELL_X8 FILLER_44_1005 ();
 FILLCELL_X4 FILLER_44_1018 ();
 FILLCELL_X2 FILLER_44_1022 ();
 FILLCELL_X1 FILLER_44_1027 ();
 FILLCELL_X2 FILLER_44_1048 ();
 FILLCELL_X4 FILLER_44_1056 ();
 FILLCELL_X1 FILLER_44_1060 ();
 FILLCELL_X8 FILLER_44_1069 ();
 FILLCELL_X1 FILLER_44_1077 ();
 FILLCELL_X1 FILLER_44_1085 ();
 FILLCELL_X2 FILLER_44_1094 ();
 FILLCELL_X1 FILLER_44_1111 ();
 FILLCELL_X8 FILLER_44_1128 ();
 FILLCELL_X2 FILLER_44_1141 ();
 FILLCELL_X1 FILLER_44_1143 ();
 FILLCELL_X2 FILLER_44_1152 ();
 FILLCELL_X4 FILLER_44_1158 ();
 FILLCELL_X2 FILLER_44_1162 ();
 FILLCELL_X1 FILLER_44_1164 ();
 FILLCELL_X2 FILLER_44_1173 ();
 FILLCELL_X8 FILLER_44_1195 ();
 FILLCELL_X4 FILLER_44_1203 ();
 FILLCELL_X2 FILLER_44_1207 ();
 FILLCELL_X32 FILLER_45_1 ();
 FILLCELL_X16 FILLER_45_33 ();
 FILLCELL_X1 FILLER_45_49 ();
 FILLCELL_X8 FILLER_45_85 ();
 FILLCELL_X4 FILLER_45_93 ();
 FILLCELL_X2 FILLER_45_97 ();
 FILLCELL_X1 FILLER_45_99 ();
 FILLCELL_X2 FILLER_45_107 ();
 FILLCELL_X1 FILLER_45_109 ();
 FILLCELL_X2 FILLER_45_113 ();
 FILLCELL_X1 FILLER_45_115 ();
 FILLCELL_X4 FILLER_45_126 ();
 FILLCELL_X2 FILLER_45_137 ();
 FILLCELL_X1 FILLER_45_139 ();
 FILLCELL_X4 FILLER_45_151 ();
 FILLCELL_X1 FILLER_45_155 ();
 FILLCELL_X2 FILLER_45_160 ();
 FILLCELL_X8 FILLER_45_170 ();
 FILLCELL_X4 FILLER_45_178 ();
 FILLCELL_X2 FILLER_45_193 ();
 FILLCELL_X1 FILLER_45_199 ();
 FILLCELL_X2 FILLER_45_204 ();
 FILLCELL_X1 FILLER_45_206 ();
 FILLCELL_X1 FILLER_45_213 ();
 FILLCELL_X32 FILLER_45_230 ();
 FILLCELL_X4 FILLER_45_262 ();
 FILLCELL_X1 FILLER_45_283 ();
 FILLCELL_X2 FILLER_45_287 ();
 FILLCELL_X1 FILLER_45_289 ();
 FILLCELL_X2 FILLER_45_320 ();
 FILLCELL_X1 FILLER_45_322 ();
 FILLCELL_X2 FILLER_45_350 ();
 FILLCELL_X1 FILLER_45_352 ();
 FILLCELL_X1 FILLER_45_363 ();
 FILLCELL_X8 FILLER_45_377 ();
 FILLCELL_X1 FILLER_45_385 ();
 FILLCELL_X2 FILLER_45_389 ();
 FILLCELL_X4 FILLER_45_395 ();
 FILLCELL_X4 FILLER_45_403 ();
 FILLCELL_X16 FILLER_45_443 ();
 FILLCELL_X32 FILLER_45_489 ();
 FILLCELL_X8 FILLER_45_521 ();
 FILLCELL_X4 FILLER_45_537 ();
 FILLCELL_X2 FILLER_45_541 ();
 FILLCELL_X1 FILLER_45_543 ();
 FILLCELL_X16 FILLER_45_550 ();
 FILLCELL_X8 FILLER_45_566 ();
 FILLCELL_X2 FILLER_45_574 ();
 FILLCELL_X1 FILLER_45_582 ();
 FILLCELL_X4 FILLER_45_606 ();
 FILLCELL_X2 FILLER_45_610 ();
 FILLCELL_X1 FILLER_45_612 ();
 FILLCELL_X4 FILLER_45_629 ();
 FILLCELL_X1 FILLER_45_633 ();
 FILLCELL_X8 FILLER_45_649 ();
 FILLCELL_X2 FILLER_45_657 ();
 FILLCELL_X16 FILLER_45_691 ();
 FILLCELL_X1 FILLER_45_707 ();
 FILLCELL_X4 FILLER_45_722 ();
 FILLCELL_X1 FILLER_45_726 ();
 FILLCELL_X8 FILLER_45_745 ();
 FILLCELL_X1 FILLER_45_777 ();
 FILLCELL_X2 FILLER_45_798 ();
 FILLCELL_X1 FILLER_45_800 ();
 FILLCELL_X2 FILLER_45_819 ();
 FILLCELL_X1 FILLER_45_821 ();
 FILLCELL_X2 FILLER_45_831 ();
 FILLCELL_X2 FILLER_45_845 ();
 FILLCELL_X2 FILLER_45_852 ();
 FILLCELL_X1 FILLER_45_854 ();
 FILLCELL_X4 FILLER_45_875 ();
 FILLCELL_X1 FILLER_45_879 ();
 FILLCELL_X8 FILLER_45_884 ();
 FILLCELL_X1 FILLER_45_892 ();
 FILLCELL_X2 FILLER_45_914 ();
 FILLCELL_X16 FILLER_45_943 ();
 FILLCELL_X16 FILLER_45_969 ();
 FILLCELL_X4 FILLER_45_985 ();
 FILLCELL_X2 FILLER_45_989 ();
 FILLCELL_X1 FILLER_45_991 ();
 FILLCELL_X2 FILLER_45_995 ();
 FILLCELL_X1 FILLER_45_997 ();
 FILLCELL_X2 FILLER_45_1011 ();
 FILLCELL_X2 FILLER_45_1036 ();
 FILLCELL_X8 FILLER_45_1042 ();
 FILLCELL_X4 FILLER_45_1050 ();
 FILLCELL_X2 FILLER_45_1054 ();
 FILLCELL_X1 FILLER_45_1066 ();
 FILLCELL_X1 FILLER_45_1077 ();
 FILLCELL_X16 FILLER_45_1081 ();
 FILLCELL_X1 FILLER_45_1097 ();
 FILLCELL_X2 FILLER_45_1124 ();
 FILLCELL_X2 FILLER_45_1152 ();
 FILLCELL_X1 FILLER_45_1166 ();
 FILLCELL_X16 FILLER_45_1183 ();
 FILLCELL_X8 FILLER_45_1199 ();
 FILLCELL_X2 FILLER_45_1207 ();
 FILLCELL_X32 FILLER_46_1 ();
 FILLCELL_X16 FILLER_46_33 ();
 FILLCELL_X4 FILLER_46_49 ();
 FILLCELL_X2 FILLER_46_53 ();
 FILLCELL_X8 FILLER_46_65 ();
 FILLCELL_X2 FILLER_46_73 ();
 FILLCELL_X4 FILLER_46_89 ();
 FILLCELL_X4 FILLER_46_105 ();
 FILLCELL_X2 FILLER_46_109 ();
 FILLCELL_X1 FILLER_46_119 ();
 FILLCELL_X2 FILLER_46_131 ();
 FILLCELL_X1 FILLER_46_133 ();
 FILLCELL_X1 FILLER_46_137 ();
 FILLCELL_X1 FILLER_46_148 ();
 FILLCELL_X4 FILLER_46_152 ();
 FILLCELL_X2 FILLER_46_156 ();
 FILLCELL_X2 FILLER_46_162 ();
 FILLCELL_X1 FILLER_46_164 ();
 FILLCELL_X2 FILLER_46_172 ();
 FILLCELL_X1 FILLER_46_185 ();
 FILLCELL_X2 FILLER_46_200 ();
 FILLCELL_X1 FILLER_46_202 ();
 FILLCELL_X2 FILLER_46_208 ();
 FILLCELL_X2 FILLER_46_214 ();
 FILLCELL_X1 FILLER_46_216 ();
 FILLCELL_X1 FILLER_46_221 ();
 FILLCELL_X16 FILLER_46_240 ();
 FILLCELL_X2 FILLER_46_256 ();
 FILLCELL_X4 FILLER_46_271 ();
 FILLCELL_X1 FILLER_46_275 ();
 FILLCELL_X2 FILLER_46_289 ();
 FILLCELL_X2 FILLER_46_309 ();
 FILLCELL_X1 FILLER_46_311 ();
 FILLCELL_X2 FILLER_46_319 ();
 FILLCELL_X1 FILLER_46_321 ();
 FILLCELL_X4 FILLER_46_327 ();
 FILLCELL_X16 FILLER_46_346 ();
 FILLCELL_X8 FILLER_46_362 ();
 FILLCELL_X2 FILLER_46_370 ();
 FILLCELL_X1 FILLER_46_372 ();
 FILLCELL_X2 FILLER_46_380 ();
 FILLCELL_X1 FILLER_46_382 ();
 FILLCELL_X4 FILLER_46_392 ();
 FILLCELL_X2 FILLER_46_396 ();
 FILLCELL_X1 FILLER_46_398 ();
 FILLCELL_X8 FILLER_46_437 ();
 FILLCELL_X4 FILLER_46_445 ();
 FILLCELL_X2 FILLER_46_449 ();
 FILLCELL_X1 FILLER_46_451 ();
 FILLCELL_X16 FILLER_46_459 ();
 FILLCELL_X1 FILLER_46_475 ();
 FILLCELL_X8 FILLER_46_504 ();
 FILLCELL_X2 FILLER_46_512 ();
 FILLCELL_X2 FILLER_46_517 ();
 FILLCELL_X1 FILLER_46_519 ();
 FILLCELL_X4 FILLER_46_523 ();
 FILLCELL_X1 FILLER_46_527 ();
 FILLCELL_X2 FILLER_46_541 ();
 FILLCELL_X8 FILLER_46_550 ();
 FILLCELL_X2 FILLER_46_558 ();
 FILLCELL_X1 FILLER_46_595 ();
 FILLCELL_X2 FILLER_46_609 ();
 FILLCELL_X8 FILLER_46_617 ();
 FILLCELL_X4 FILLER_46_632 ();
 FILLCELL_X2 FILLER_46_636 ();
 FILLCELL_X1 FILLER_46_638 ();
 FILLCELL_X2 FILLER_46_659 ();
 FILLCELL_X4 FILLER_46_702 ();
 FILLCELL_X2 FILLER_46_706 ();
 FILLCELL_X1 FILLER_46_708 ();
 FILLCELL_X8 FILLER_46_721 ();
 FILLCELL_X4 FILLER_46_729 ();
 FILLCELL_X2 FILLER_46_733 ();
 FILLCELL_X1 FILLER_46_735 ();
 FILLCELL_X1 FILLER_46_762 ();
 FILLCELL_X4 FILLER_46_783 ();
 FILLCELL_X2 FILLER_46_787 ();
 FILLCELL_X1 FILLER_46_789 ();
 FILLCELL_X2 FILLER_46_797 ();
 FILLCELL_X1 FILLER_46_799 ();
 FILLCELL_X2 FILLER_46_804 ();
 FILLCELL_X8 FILLER_46_822 ();
 FILLCELL_X2 FILLER_46_838 ();
 FILLCELL_X8 FILLER_46_844 ();
 FILLCELL_X2 FILLER_46_852 ();
 FILLCELL_X1 FILLER_46_854 ();
 FILLCELL_X8 FILLER_46_875 ();
 FILLCELL_X1 FILLER_46_883 ();
 FILLCELL_X8 FILLER_46_895 ();
 FILLCELL_X1 FILLER_46_903 ();
 FILLCELL_X2 FILLER_46_907 ();
 FILLCELL_X4 FILLER_46_916 ();
 FILLCELL_X8 FILLER_46_932 ();
 FILLCELL_X4 FILLER_46_940 ();
 FILLCELL_X2 FILLER_46_944 ();
 FILLCELL_X1 FILLER_46_946 ();
 FILLCELL_X4 FILLER_46_954 ();
 FILLCELL_X32 FILLER_46_971 ();
 FILLCELL_X4 FILLER_46_1003 ();
 FILLCELL_X2 FILLER_46_1007 ();
 FILLCELL_X1 FILLER_46_1009 ();
 FILLCELL_X2 FILLER_46_1030 ();
 FILLCELL_X1 FILLER_46_1032 ();
 FILLCELL_X4 FILLER_46_1039 ();
 FILLCELL_X1 FILLER_46_1043 ();
 FILLCELL_X1 FILLER_46_1049 ();
 FILLCELL_X4 FILLER_46_1061 ();
 FILLCELL_X2 FILLER_46_1065 ();
 FILLCELL_X16 FILLER_46_1086 ();
 FILLCELL_X8 FILLER_46_1102 ();
 FILLCELL_X4 FILLER_46_1110 ();
 FILLCELL_X1 FILLER_46_1114 ();
 FILLCELL_X2 FILLER_46_1118 ();
 FILLCELL_X2 FILLER_46_1123 ();
 FILLCELL_X2 FILLER_46_1129 ();
 FILLCELL_X2 FILLER_46_1135 ();
 FILLCELL_X1 FILLER_46_1137 ();
 FILLCELL_X1 FILLER_46_1144 ();
 FILLCELL_X2 FILLER_46_1152 ();
 FILLCELL_X1 FILLER_46_1154 ();
 FILLCELL_X4 FILLER_46_1163 ();
 FILLCELL_X2 FILLER_46_1167 ();
 FILLCELL_X1 FILLER_46_1169 ();
 FILLCELL_X4 FILLER_46_1200 ();
 FILLCELL_X1 FILLER_46_1204 ();
 FILLCELL_X32 FILLER_47_1 ();
 FILLCELL_X16 FILLER_47_33 ();
 FILLCELL_X2 FILLER_47_49 ();
 FILLCELL_X1 FILLER_47_61 ();
 FILLCELL_X1 FILLER_47_73 ();
 FILLCELL_X4 FILLER_47_78 ();
 FILLCELL_X2 FILLER_47_82 ();
 FILLCELL_X1 FILLER_47_84 ();
 FILLCELL_X4 FILLER_47_111 ();
 FILLCELL_X2 FILLER_47_115 ();
 FILLCELL_X1 FILLER_47_117 ();
 FILLCELL_X8 FILLER_47_122 ();
 FILLCELL_X1 FILLER_47_135 ();
 FILLCELL_X1 FILLER_47_141 ();
 FILLCELL_X1 FILLER_47_152 ();
 FILLCELL_X2 FILLER_47_193 ();
 FILLCELL_X1 FILLER_47_195 ();
 FILLCELL_X8 FILLER_47_200 ();
 FILLCELL_X32 FILLER_47_222 ();
 FILLCELL_X4 FILLER_47_254 ();
 FILLCELL_X1 FILLER_47_258 ();
 FILLCELL_X4 FILLER_47_272 ();
 FILLCELL_X2 FILLER_47_276 ();
 FILLCELL_X16 FILLER_47_334 ();
 FILLCELL_X1 FILLER_47_350 ();
 FILLCELL_X1 FILLER_47_358 ();
 FILLCELL_X2 FILLER_47_366 ();
 FILLCELL_X2 FILLER_47_379 ();
 FILLCELL_X1 FILLER_47_381 ();
 FILLCELL_X1 FILLER_47_409 ();
 FILLCELL_X2 FILLER_47_418 ();
 FILLCELL_X2 FILLER_47_428 ();
 FILLCELL_X1 FILLER_47_430 ();
 FILLCELL_X16 FILLER_47_435 ();
 FILLCELL_X4 FILLER_47_451 ();
 FILLCELL_X2 FILLER_47_455 ();
 FILLCELL_X1 FILLER_47_457 ();
 FILLCELL_X8 FILLER_47_471 ();
 FILLCELL_X2 FILLER_47_479 ();
 FILLCELL_X1 FILLER_47_481 ();
 FILLCELL_X2 FILLER_47_486 ();
 FILLCELL_X1 FILLER_47_488 ();
 FILLCELL_X2 FILLER_47_495 ();
 FILLCELL_X1 FILLER_47_497 ();
 FILLCELL_X1 FILLER_47_522 ();
 FILLCELL_X2 FILLER_47_554 ();
 FILLCELL_X1 FILLER_47_556 ();
 FILLCELL_X1 FILLER_47_576 ();
 FILLCELL_X1 FILLER_47_586 ();
 FILLCELL_X1 FILLER_47_630 ();
 FILLCELL_X1 FILLER_47_635 ();
 FILLCELL_X1 FILLER_47_646 ();
 FILLCELL_X2 FILLER_47_652 ();
 FILLCELL_X1 FILLER_47_663 ();
 FILLCELL_X8 FILLER_47_674 ();
 FILLCELL_X4 FILLER_47_682 ();
 FILLCELL_X32 FILLER_47_691 ();
 FILLCELL_X32 FILLER_47_723 ();
 FILLCELL_X1 FILLER_47_755 ();
 FILLCELL_X4 FILLER_47_769 ();
 FILLCELL_X4 FILLER_47_793 ();
 FILLCELL_X2 FILLER_47_814 ();
 FILLCELL_X4 FILLER_47_852 ();
 FILLCELL_X4 FILLER_47_865 ();
 FILLCELL_X4 FILLER_47_873 ();
 FILLCELL_X1 FILLER_47_877 ();
 FILLCELL_X1 FILLER_47_889 ();
 FILLCELL_X8 FILLER_47_910 ();
 FILLCELL_X4 FILLER_47_918 ();
 FILLCELL_X1 FILLER_47_922 ();
 FILLCELL_X8 FILLER_47_930 ();
 FILLCELL_X1 FILLER_47_938 ();
 FILLCELL_X4 FILLER_47_953 ();
 FILLCELL_X2 FILLER_47_957 ();
 FILLCELL_X1 FILLER_47_959 ();
 FILLCELL_X16 FILLER_47_993 ();
 FILLCELL_X8 FILLER_47_1009 ();
 FILLCELL_X1 FILLER_47_1017 ();
 FILLCELL_X4 FILLER_47_1025 ();
 FILLCELL_X1 FILLER_47_1044 ();
 FILLCELL_X1 FILLER_47_1051 ();
 FILLCELL_X4 FILLER_47_1058 ();
 FILLCELL_X1 FILLER_47_1062 ();
 FILLCELL_X4 FILLER_47_1066 ();
 FILLCELL_X2 FILLER_47_1070 ();
 FILLCELL_X8 FILLER_47_1091 ();
 FILLCELL_X8 FILLER_47_1118 ();
 FILLCELL_X2 FILLER_47_1150 ();
 FILLCELL_X1 FILLER_47_1152 ();
 FILLCELL_X1 FILLER_47_1157 ();
 FILLCELL_X1 FILLER_47_1173 ();
 FILLCELL_X8 FILLER_47_1181 ();
 FILLCELL_X2 FILLER_47_1189 ();
 FILLCELL_X8 FILLER_47_1194 ();
 FILLCELL_X4 FILLER_47_1202 ();
 FILLCELL_X2 FILLER_47_1206 ();
 FILLCELL_X1 FILLER_47_1208 ();
 FILLCELL_X32 FILLER_48_1 ();
 FILLCELL_X32 FILLER_48_33 ();
 FILLCELL_X2 FILLER_48_65 ();
 FILLCELL_X2 FILLER_48_71 ();
 FILLCELL_X1 FILLER_48_73 ();
 FILLCELL_X2 FILLER_48_78 ();
 FILLCELL_X2 FILLER_48_103 ();
 FILLCELL_X1 FILLER_48_105 ();
 FILLCELL_X1 FILLER_48_117 ();
 FILLCELL_X1 FILLER_48_122 ();
 FILLCELL_X2 FILLER_48_137 ();
 FILLCELL_X4 FILLER_48_168 ();
 FILLCELL_X2 FILLER_48_172 ();
 FILLCELL_X1 FILLER_48_174 ();
 FILLCELL_X8 FILLER_48_178 ();
 FILLCELL_X4 FILLER_48_186 ();
 FILLCELL_X2 FILLER_48_190 ();
 FILLCELL_X2 FILLER_48_196 ();
 FILLCELL_X4 FILLER_48_204 ();
 FILLCELL_X4 FILLER_48_212 ();
 FILLCELL_X2 FILLER_48_225 ();
 FILLCELL_X16 FILLER_48_240 ();
 FILLCELL_X4 FILLER_48_256 ();
 FILLCELL_X2 FILLER_48_260 ();
 FILLCELL_X1 FILLER_48_262 ();
 FILLCELL_X1 FILLER_48_268 ();
 FILLCELL_X2 FILLER_48_282 ();
 FILLCELL_X1 FILLER_48_325 ();
 FILLCELL_X4 FILLER_48_344 ();
 FILLCELL_X2 FILLER_48_348 ();
 FILLCELL_X4 FILLER_48_361 ();
 FILLCELL_X2 FILLER_48_365 ();
 FILLCELL_X2 FILLER_48_385 ();
 FILLCELL_X1 FILLER_48_387 ();
 FILLCELL_X1 FILLER_48_401 ();
 FILLCELL_X2 FILLER_48_406 ();
 FILLCELL_X1 FILLER_48_408 ();
 FILLCELL_X2 FILLER_48_415 ();
 FILLCELL_X1 FILLER_48_417 ();
 FILLCELL_X8 FILLER_48_439 ();
 FILLCELL_X4 FILLER_48_447 ();
 FILLCELL_X2 FILLER_48_451 ();
 FILLCELL_X16 FILLER_48_462 ();
 FILLCELL_X8 FILLER_48_478 ();
 FILLCELL_X2 FILLER_48_486 ();
 FILLCELL_X1 FILLER_48_488 ();
 FILLCELL_X4 FILLER_48_506 ();
 FILLCELL_X1 FILLER_48_510 ();
 FILLCELL_X2 FILLER_48_534 ();
 FILLCELL_X4 FILLER_48_567 ();
 FILLCELL_X1 FILLER_48_571 ();
 FILLCELL_X8 FILLER_48_594 ();
 FILLCELL_X2 FILLER_48_616 ();
 FILLCELL_X1 FILLER_48_618 ();
 FILLCELL_X8 FILLER_48_622 ();
 FILLCELL_X1 FILLER_48_630 ();
 FILLCELL_X1 FILLER_48_673 ();
 FILLCELL_X4 FILLER_48_691 ();
 FILLCELL_X1 FILLER_48_695 ();
 FILLCELL_X32 FILLER_48_709 ();
 FILLCELL_X2 FILLER_48_741 ();
 FILLCELL_X1 FILLER_48_743 ();
 FILLCELL_X4 FILLER_48_764 ();
 FILLCELL_X2 FILLER_48_768 ();
 FILLCELL_X2 FILLER_48_783 ();
 FILLCELL_X1 FILLER_48_805 ();
 FILLCELL_X2 FILLER_48_824 ();
 FILLCELL_X1 FILLER_48_826 ();
 FILLCELL_X2 FILLER_48_834 ();
 FILLCELL_X1 FILLER_48_836 ();
 FILLCELL_X2 FILLER_48_852 ();
 FILLCELL_X1 FILLER_48_854 ();
 FILLCELL_X2 FILLER_48_858 ();
 FILLCELL_X8 FILLER_48_895 ();
 FILLCELL_X2 FILLER_48_903 ();
 FILLCELL_X1 FILLER_48_905 ();
 FILLCELL_X32 FILLER_48_919 ();
 FILLCELL_X32 FILLER_48_951 ();
 FILLCELL_X16 FILLER_48_983 ();
 FILLCELL_X8 FILLER_48_999 ();
 FILLCELL_X2 FILLER_48_1007 ();
 FILLCELL_X1 FILLER_48_1009 ();
 FILLCELL_X4 FILLER_48_1037 ();
 FILLCELL_X1 FILLER_48_1041 ();
 FILLCELL_X8 FILLER_48_1056 ();
 FILLCELL_X4 FILLER_48_1086 ();
 FILLCELL_X1 FILLER_48_1107 ();
 FILLCELL_X1 FILLER_48_1115 ();
 FILLCELL_X4 FILLER_48_1139 ();
 FILLCELL_X2 FILLER_48_1143 ();
 FILLCELL_X1 FILLER_48_1145 ();
 FILLCELL_X4 FILLER_48_1149 ();
 FILLCELL_X2 FILLER_48_1157 ();
 FILLCELL_X1 FILLER_48_1159 ();
 FILLCELL_X8 FILLER_48_1165 ();
 FILLCELL_X4 FILLER_48_1173 ();
 FILLCELL_X2 FILLER_48_1177 ();
 FILLCELL_X4 FILLER_48_1194 ();
 FILLCELL_X1 FILLER_48_1198 ();
 FILLCELL_X2 FILLER_48_1202 ();
 FILLCELL_X1 FILLER_48_1204 ();
 FILLCELL_X1 FILLER_48_1208 ();
 FILLCELL_X32 FILLER_49_1 ();
 FILLCELL_X16 FILLER_49_33 ();
 FILLCELL_X8 FILLER_49_49 ();
 FILLCELL_X2 FILLER_49_82 ();
 FILLCELL_X2 FILLER_49_91 ();
 FILLCELL_X2 FILLER_49_100 ();
 FILLCELL_X1 FILLER_49_112 ();
 FILLCELL_X2 FILLER_49_117 ();
 FILLCELL_X2 FILLER_49_124 ();
 FILLCELL_X2 FILLER_49_129 ();
 FILLCELL_X2 FILLER_49_134 ();
 FILLCELL_X1 FILLER_49_136 ();
 FILLCELL_X2 FILLER_49_148 ();
 FILLCELL_X4 FILLER_49_153 ();
 FILLCELL_X1 FILLER_49_157 ();
 FILLCELL_X2 FILLER_49_165 ();
 FILLCELL_X1 FILLER_49_167 ();
 FILLCELL_X4 FILLER_49_177 ();
 FILLCELL_X4 FILLER_49_186 ();
 FILLCELL_X2 FILLER_49_190 ();
 FILLCELL_X1 FILLER_49_202 ();
 FILLCELL_X1 FILLER_49_214 ();
 FILLCELL_X32 FILLER_49_223 ();
 FILLCELL_X4 FILLER_49_255 ();
 FILLCELL_X8 FILLER_49_272 ();
 FILLCELL_X1 FILLER_49_280 ();
 FILLCELL_X2 FILLER_49_297 ();
 FILLCELL_X1 FILLER_49_299 ();
 FILLCELL_X1 FILLER_49_311 ();
 FILLCELL_X1 FILLER_49_326 ();
 FILLCELL_X8 FILLER_49_334 ();
 FILLCELL_X4 FILLER_49_342 ();
 FILLCELL_X2 FILLER_49_351 ();
 FILLCELL_X4 FILLER_49_378 ();
 FILLCELL_X2 FILLER_49_382 ();
 FILLCELL_X1 FILLER_49_384 ();
 FILLCELL_X2 FILLER_49_393 ();
 FILLCELL_X2 FILLER_49_399 ();
 FILLCELL_X2 FILLER_49_405 ();
 FILLCELL_X1 FILLER_49_407 ();
 FILLCELL_X2 FILLER_49_412 ();
 FILLCELL_X1 FILLER_49_414 ();
 FILLCELL_X16 FILLER_49_429 ();
 FILLCELL_X4 FILLER_49_445 ();
 FILLCELL_X2 FILLER_49_449 ();
 FILLCELL_X1 FILLER_49_451 ();
 FILLCELL_X32 FILLER_49_492 ();
 FILLCELL_X2 FILLER_49_524 ();
 FILLCELL_X1 FILLER_49_526 ();
 FILLCELL_X2 FILLER_49_533 ();
 FILLCELL_X1 FILLER_49_535 ();
 FILLCELL_X8 FILLER_49_563 ();
 FILLCELL_X2 FILLER_49_593 ();
 FILLCELL_X1 FILLER_49_595 ();
 FILLCELL_X2 FILLER_49_606 ();
 FILLCELL_X1 FILLER_49_608 ();
 FILLCELL_X2 FILLER_49_622 ();
 FILLCELL_X2 FILLER_49_633 ();
 FILLCELL_X8 FILLER_49_645 ();
 FILLCELL_X2 FILLER_49_653 ();
 FILLCELL_X1 FILLER_49_655 ();
 FILLCELL_X16 FILLER_49_661 ();
 FILLCELL_X8 FILLER_49_677 ();
 FILLCELL_X1 FILLER_49_685 ();
 FILLCELL_X8 FILLER_49_690 ();
 FILLCELL_X4 FILLER_49_698 ();
 FILLCELL_X2 FILLER_49_702 ();
 FILLCELL_X1 FILLER_49_704 ();
 FILLCELL_X32 FILLER_49_722 ();
 FILLCELL_X32 FILLER_49_754 ();
 FILLCELL_X16 FILLER_49_786 ();
 FILLCELL_X4 FILLER_49_802 ();
 FILLCELL_X1 FILLER_49_806 ();
 FILLCELL_X8 FILLER_49_820 ();
 FILLCELL_X4 FILLER_49_828 ();
 FILLCELL_X4 FILLER_49_843 ();
 FILLCELL_X1 FILLER_49_847 ();
 FILLCELL_X8 FILLER_49_877 ();
 FILLCELL_X4 FILLER_49_885 ();
 FILLCELL_X1 FILLER_49_889 ();
 FILLCELL_X4 FILLER_49_894 ();
 FILLCELL_X2 FILLER_49_902 ();
 FILLCELL_X4 FILLER_49_913 ();
 FILLCELL_X16 FILLER_49_921 ();
 FILLCELL_X1 FILLER_49_937 ();
 FILLCELL_X8 FILLER_49_968 ();
 FILLCELL_X1 FILLER_49_976 ();
 FILLCELL_X16 FILLER_49_996 ();
 FILLCELL_X4 FILLER_49_1012 ();
 FILLCELL_X2 FILLER_49_1016 ();
 FILLCELL_X1 FILLER_49_1018 ();
 FILLCELL_X1 FILLER_49_1024 ();
 FILLCELL_X4 FILLER_49_1046 ();
 FILLCELL_X4 FILLER_49_1061 ();
 FILLCELL_X2 FILLER_49_1077 ();
 FILLCELL_X4 FILLER_49_1098 ();
 FILLCELL_X4 FILLER_49_1111 ();
 FILLCELL_X2 FILLER_49_1115 ();
 FILLCELL_X4 FILLER_49_1120 ();
 FILLCELL_X2 FILLER_49_1124 ();
 FILLCELL_X1 FILLER_49_1126 ();
 FILLCELL_X2 FILLER_49_1133 ();
 FILLCELL_X8 FILLER_49_1155 ();
 FILLCELL_X4 FILLER_49_1166 ();
 FILLCELL_X2 FILLER_49_1170 ();
 FILLCELL_X16 FILLER_49_1182 ();
 FILLCELL_X8 FILLER_49_1198 ();
 FILLCELL_X2 FILLER_49_1206 ();
 FILLCELL_X1 FILLER_49_1208 ();
 FILLCELL_X32 FILLER_50_1 ();
 FILLCELL_X8 FILLER_50_33 ();
 FILLCELL_X4 FILLER_50_41 ();
 FILLCELL_X2 FILLER_50_45 ();
 FILLCELL_X1 FILLER_50_99 ();
 FILLCELL_X1 FILLER_50_111 ();
 FILLCELL_X2 FILLER_50_124 ();
 FILLCELL_X1 FILLER_50_126 ();
 FILLCELL_X1 FILLER_50_135 ();
 FILLCELL_X1 FILLER_50_143 ();
 FILLCELL_X4 FILLER_50_157 ();
 FILLCELL_X4 FILLER_50_164 ();
 FILLCELL_X1 FILLER_50_168 ();
 FILLCELL_X4 FILLER_50_174 ();
 FILLCELL_X1 FILLER_50_178 ();
 FILLCELL_X4 FILLER_50_184 ();
 FILLCELL_X2 FILLER_50_188 ();
 FILLCELL_X1 FILLER_50_190 ();
 FILLCELL_X2 FILLER_50_201 ();
 FILLCELL_X4 FILLER_50_214 ();
 FILLCELL_X1 FILLER_50_218 ();
 FILLCELL_X16 FILLER_50_226 ();
 FILLCELL_X8 FILLER_50_242 ();
 FILLCELL_X2 FILLER_50_250 ();
 FILLCELL_X4 FILLER_50_271 ();
 FILLCELL_X1 FILLER_50_275 ();
 FILLCELL_X1 FILLER_50_287 ();
 FILLCELL_X1 FILLER_50_291 ();
 FILLCELL_X8 FILLER_50_337 ();
 FILLCELL_X2 FILLER_50_345 ();
 FILLCELL_X1 FILLER_50_347 ();
 FILLCELL_X2 FILLER_50_360 ();
 FILLCELL_X1 FILLER_50_362 ();
 FILLCELL_X2 FILLER_50_367 ();
 FILLCELL_X1 FILLER_50_369 ();
 FILLCELL_X8 FILLER_50_377 ();
 FILLCELL_X8 FILLER_50_389 ();
 FILLCELL_X4 FILLER_50_397 ();
 FILLCELL_X2 FILLER_50_401 ();
 FILLCELL_X32 FILLER_50_427 ();
 FILLCELL_X16 FILLER_50_459 ();
 FILLCELL_X1 FILLER_50_490 ();
 FILLCELL_X2 FILLER_50_494 ();
 FILLCELL_X1 FILLER_50_496 ();
 FILLCELL_X8 FILLER_50_525 ();
 FILLCELL_X4 FILLER_50_533 ();
 FILLCELL_X2 FILLER_50_537 ();
 FILLCELL_X1 FILLER_50_539 ();
 FILLCELL_X16 FILLER_50_570 ();
 FILLCELL_X8 FILLER_50_586 ();
 FILLCELL_X1 FILLER_50_610 ();
 FILLCELL_X16 FILLER_50_654 ();
 FILLCELL_X8 FILLER_50_670 ();
 FILLCELL_X4 FILLER_50_678 ();
 FILLCELL_X1 FILLER_50_682 ();
 FILLCELL_X4 FILLER_50_700 ();
 FILLCELL_X1 FILLER_50_704 ();
 FILLCELL_X32 FILLER_50_712 ();
 FILLCELL_X32 FILLER_50_744 ();
 FILLCELL_X4 FILLER_50_776 ();
 FILLCELL_X2 FILLER_50_780 ();
 FILLCELL_X1 FILLER_50_782 ();
 FILLCELL_X16 FILLER_50_800 ();
 FILLCELL_X8 FILLER_50_816 ();
 FILLCELL_X1 FILLER_50_824 ();
 FILLCELL_X2 FILLER_50_838 ();
 FILLCELL_X1 FILLER_50_840 ();
 FILLCELL_X4 FILLER_50_845 ();
 FILLCELL_X2 FILLER_50_849 ();
 FILLCELL_X4 FILLER_50_862 ();
 FILLCELL_X2 FILLER_50_866 ();
 FILLCELL_X1 FILLER_50_872 ();
 FILLCELL_X1 FILLER_50_877 ();
 FILLCELL_X1 FILLER_50_886 ();
 FILLCELL_X1 FILLER_50_891 ();
 FILLCELL_X1 FILLER_50_896 ();
 FILLCELL_X1 FILLER_50_901 ();
 FILLCELL_X32 FILLER_50_906 ();
 FILLCELL_X4 FILLER_50_962 ();
 FILLCELL_X2 FILLER_50_966 ();
 FILLCELL_X1 FILLER_50_968 ();
 FILLCELL_X2 FILLER_50_989 ();
 FILLCELL_X1 FILLER_50_991 ();
 FILLCELL_X8 FILLER_50_1011 ();
 FILLCELL_X1 FILLER_50_1019 ();
 FILLCELL_X4 FILLER_50_1048 ();
 FILLCELL_X2 FILLER_50_1052 ();
 FILLCELL_X1 FILLER_50_1054 ();
 FILLCELL_X8 FILLER_50_1062 ();
 FILLCELL_X2 FILLER_50_1070 ();
 FILLCELL_X4 FILLER_50_1080 ();
 FILLCELL_X8 FILLER_50_1092 ();
 FILLCELL_X2 FILLER_50_1100 ();
 FILLCELL_X1 FILLER_50_1102 ();
 FILLCELL_X1 FILLER_50_1113 ();
 FILLCELL_X1 FILLER_50_1129 ();
 FILLCELL_X1 FILLER_50_1140 ();
 FILLCELL_X4 FILLER_50_1153 ();
 FILLCELL_X1 FILLER_50_1157 ();
 FILLCELL_X1 FILLER_50_1165 ();
 FILLCELL_X2 FILLER_50_1176 ();
 FILLCELL_X1 FILLER_50_1178 ();
 FILLCELL_X2 FILLER_50_1187 ();
 FILLCELL_X16 FILLER_50_1192 ();
 FILLCELL_X1 FILLER_50_1208 ();
 FILLCELL_X16 FILLER_51_1 ();
 FILLCELL_X8 FILLER_51_17 ();
 FILLCELL_X4 FILLER_51_25 ();
 FILLCELL_X2 FILLER_51_29 ();
 FILLCELL_X32 FILLER_51_34 ();
 FILLCELL_X1 FILLER_51_66 ();
 FILLCELL_X2 FILLER_51_95 ();
 FILLCELL_X2 FILLER_51_110 ();
 FILLCELL_X1 FILLER_51_112 ();
 FILLCELL_X4 FILLER_51_120 ();
 FILLCELL_X2 FILLER_51_124 ();
 FILLCELL_X1 FILLER_51_132 ();
 FILLCELL_X2 FILLER_51_163 ();
 FILLCELL_X1 FILLER_51_171 ();
 FILLCELL_X2 FILLER_51_175 ();
 FILLCELL_X1 FILLER_51_177 ();
 FILLCELL_X2 FILLER_51_200 ();
 FILLCELL_X32 FILLER_51_209 ();
 FILLCELL_X16 FILLER_51_241 ();
 FILLCELL_X1 FILLER_51_257 ();
 FILLCELL_X4 FILLER_51_272 ();
 FILLCELL_X2 FILLER_51_276 ();
 FILLCELL_X1 FILLER_51_311 ();
 FILLCELL_X2 FILLER_51_325 ();
 FILLCELL_X1 FILLER_51_342 ();
 FILLCELL_X1 FILLER_51_346 ();
 FILLCELL_X2 FILLER_51_354 ();
 FILLCELL_X1 FILLER_51_356 ();
 FILLCELL_X1 FILLER_51_367 ();
 FILLCELL_X1 FILLER_51_372 ();
 FILLCELL_X2 FILLER_51_384 ();
 FILLCELL_X1 FILLER_51_386 ();
 FILLCELL_X8 FILLER_51_391 ();
 FILLCELL_X4 FILLER_51_399 ();
 FILLCELL_X2 FILLER_51_403 ();
 FILLCELL_X1 FILLER_51_405 ();
 FILLCELL_X8 FILLER_51_424 ();
 FILLCELL_X4 FILLER_51_432 ();
 FILLCELL_X2 FILLER_51_436 ();
 FILLCELL_X1 FILLER_51_438 ();
 FILLCELL_X2 FILLER_51_456 ();
 FILLCELL_X1 FILLER_51_458 ();
 FILLCELL_X2 FILLER_51_472 ();
 FILLCELL_X1 FILLER_51_520 ();
 FILLCELL_X4 FILLER_51_528 ();
 FILLCELL_X2 FILLER_51_532 ();
 FILLCELL_X16 FILLER_51_540 ();
 FILLCELL_X4 FILLER_51_556 ();
 FILLCELL_X2 FILLER_51_560 ();
 FILLCELL_X1 FILLER_51_562 ();
 FILLCELL_X1 FILLER_51_576 ();
 FILLCELL_X2 FILLER_51_588 ();
 FILLCELL_X1 FILLER_51_590 ();
 FILLCELL_X2 FILLER_51_628 ();
 FILLCELL_X1 FILLER_51_653 ();
 FILLCELL_X8 FILLER_51_682 ();
 FILLCELL_X2 FILLER_51_690 ();
 FILLCELL_X1 FILLER_51_692 ();
 FILLCELL_X8 FILLER_51_722 ();
 FILLCELL_X4 FILLER_51_730 ();
 FILLCELL_X2 FILLER_51_734 ();
 FILLCELL_X1 FILLER_51_736 ();
 FILLCELL_X2 FILLER_51_747 ();
 FILLCELL_X16 FILLER_51_753 ();
 FILLCELL_X4 FILLER_51_769 ();
 FILLCELL_X2 FILLER_51_773 ();
 FILLCELL_X8 FILLER_51_779 ();
 FILLCELL_X2 FILLER_51_787 ();
 FILLCELL_X1 FILLER_51_789 ();
 FILLCELL_X16 FILLER_51_795 ();
 FILLCELL_X4 FILLER_51_811 ();
 FILLCELL_X1 FILLER_51_815 ();
 FILLCELL_X16 FILLER_51_823 ();
 FILLCELL_X1 FILLER_51_839 ();
 FILLCELL_X8 FILLER_51_878 ();
 FILLCELL_X16 FILLER_51_893 ();
 FILLCELL_X8 FILLER_51_928 ();
 FILLCELL_X4 FILLER_51_936 ();
 FILLCELL_X8 FILLER_51_946 ();
 FILLCELL_X2 FILLER_51_967 ();
 FILLCELL_X1 FILLER_51_969 ();
 FILLCELL_X16 FILLER_51_1002 ();
 FILLCELL_X4 FILLER_51_1018 ();
 FILLCELL_X2 FILLER_51_1022 ();
 FILLCELL_X8 FILLER_51_1031 ();
 FILLCELL_X2 FILLER_51_1039 ();
 FILLCELL_X2 FILLER_51_1048 ();
 FILLCELL_X1 FILLER_51_1050 ();
 FILLCELL_X4 FILLER_51_1054 ();
 FILLCELL_X1 FILLER_51_1069 ();
 FILLCELL_X2 FILLER_51_1073 ();
 FILLCELL_X1 FILLER_51_1075 ();
 FILLCELL_X4 FILLER_51_1091 ();
 FILLCELL_X2 FILLER_51_1134 ();
 FILLCELL_X1 FILLER_51_1136 ();
 FILLCELL_X2 FILLER_51_1155 ();
 FILLCELL_X8 FILLER_51_1177 ();
 FILLCELL_X2 FILLER_51_1185 ();
 FILLCELL_X1 FILLER_51_1187 ();
 FILLCELL_X16 FILLER_51_1191 ();
 FILLCELL_X2 FILLER_51_1207 ();
 FILLCELL_X32 FILLER_52_1 ();
 FILLCELL_X4 FILLER_52_33 ();
 FILLCELL_X1 FILLER_52_37 ();
 FILLCELL_X4 FILLER_52_53 ();
 FILLCELL_X1 FILLER_52_57 ();
 FILLCELL_X2 FILLER_52_73 ();
 FILLCELL_X1 FILLER_52_75 ();
 FILLCELL_X2 FILLER_52_90 ();
 FILLCELL_X1 FILLER_52_92 ();
 FILLCELL_X2 FILLER_52_98 ();
 FILLCELL_X1 FILLER_52_100 ();
 FILLCELL_X2 FILLER_52_110 ();
 FILLCELL_X1 FILLER_52_112 ();
 FILLCELL_X4 FILLER_52_132 ();
 FILLCELL_X1 FILLER_52_136 ();
 FILLCELL_X1 FILLER_52_147 ();
 FILLCELL_X2 FILLER_52_153 ();
 FILLCELL_X2 FILLER_52_173 ();
 FILLCELL_X1 FILLER_52_195 ();
 FILLCELL_X8 FILLER_52_200 ();
 FILLCELL_X32 FILLER_52_213 ();
 FILLCELL_X4 FILLER_52_245 ();
 FILLCELL_X1 FILLER_52_249 ();
 FILLCELL_X4 FILLER_52_264 ();
 FILLCELL_X2 FILLER_52_268 ();
 FILLCELL_X1 FILLER_52_270 ();
 FILLCELL_X1 FILLER_52_278 ();
 FILLCELL_X1 FILLER_52_286 ();
 FILLCELL_X2 FILLER_52_313 ();
 FILLCELL_X4 FILLER_52_322 ();
 FILLCELL_X2 FILLER_52_326 ();
 FILLCELL_X8 FILLER_52_337 ();
 FILLCELL_X8 FILLER_52_353 ();
 FILLCELL_X4 FILLER_52_361 ();
 FILLCELL_X4 FILLER_52_369 ();
 FILLCELL_X2 FILLER_52_373 ();
 FILLCELL_X4 FILLER_52_399 ();
 FILLCELL_X1 FILLER_52_406 ();
 FILLCELL_X16 FILLER_52_429 ();
 FILLCELL_X8 FILLER_52_445 ();
 FILLCELL_X2 FILLER_52_453 ();
 FILLCELL_X1 FILLER_52_455 ();
 FILLCELL_X4 FILLER_52_461 ();
 FILLCELL_X1 FILLER_52_465 ();
 FILLCELL_X1 FILLER_52_479 ();
 FILLCELL_X4 FILLER_52_482 ();
 FILLCELL_X2 FILLER_52_486 ();
 FILLCELL_X1 FILLER_52_488 ();
 FILLCELL_X16 FILLER_52_513 ();
 FILLCELL_X1 FILLER_52_529 ();
 FILLCELL_X2 FILLER_52_537 ();
 FILLCELL_X1 FILLER_52_539 ();
 FILLCELL_X2 FILLER_52_544 ();
 FILLCELL_X1 FILLER_52_602 ();
 FILLCELL_X1 FILLER_52_609 ();
 FILLCELL_X1 FILLER_52_626 ();
 FILLCELL_X1 FILLER_52_630 ();
 FILLCELL_X16 FILLER_52_655 ();
 FILLCELL_X4 FILLER_52_671 ();
 FILLCELL_X1 FILLER_52_678 ();
 FILLCELL_X16 FILLER_52_683 ();
 FILLCELL_X4 FILLER_52_699 ();
 FILLCELL_X2 FILLER_52_703 ();
 FILLCELL_X16 FILLER_52_709 ();
 FILLCELL_X8 FILLER_52_725 ();
 FILLCELL_X4 FILLER_52_733 ();
 FILLCELL_X32 FILLER_52_740 ();
 FILLCELL_X4 FILLER_52_772 ();
 FILLCELL_X2 FILLER_52_793 ();
 FILLCELL_X1 FILLER_52_795 ();
 FILLCELL_X32 FILLER_52_803 ();
 FILLCELL_X32 FILLER_52_835 ();
 FILLCELL_X16 FILLER_52_867 ();
 FILLCELL_X8 FILLER_52_883 ();
 FILLCELL_X4 FILLER_52_891 ();
 FILLCELL_X16 FILLER_52_912 ();
 FILLCELL_X4 FILLER_52_928 ();
 FILLCELL_X2 FILLER_52_932 ();
 FILLCELL_X1 FILLER_52_934 ();
 FILLCELL_X1 FILLER_52_957 ();
 FILLCELL_X1 FILLER_52_964 ();
 FILLCELL_X1 FILLER_52_971 ();
 FILLCELL_X4 FILLER_52_978 ();
 FILLCELL_X2 FILLER_52_982 ();
 FILLCELL_X1 FILLER_52_984 ();
 FILLCELL_X16 FILLER_52_1002 ();
 FILLCELL_X2 FILLER_52_1018 ();
 FILLCELL_X1 FILLER_52_1027 ();
 FILLCELL_X4 FILLER_52_1035 ();
 FILLCELL_X4 FILLER_52_1047 ();
 FILLCELL_X1 FILLER_52_1057 ();
 FILLCELL_X1 FILLER_52_1061 ();
 FILLCELL_X1 FILLER_52_1072 ();
 FILLCELL_X8 FILLER_52_1084 ();
 FILLCELL_X1 FILLER_52_1096 ();
 FILLCELL_X8 FILLER_52_1115 ();
 FILLCELL_X1 FILLER_52_1123 ();
 FILLCELL_X1 FILLER_52_1128 ();
 FILLCELL_X2 FILLER_52_1133 ();
 FILLCELL_X1 FILLER_52_1135 ();
 FILLCELL_X8 FILLER_52_1139 ();
 FILLCELL_X4 FILLER_52_1147 ();
 FILLCELL_X4 FILLER_52_1155 ();
 FILLCELL_X8 FILLER_52_1163 ();
 FILLCELL_X2 FILLER_52_1171 ();
 FILLCELL_X2 FILLER_52_1177 ();
 FILLCELL_X1 FILLER_52_1179 ();
 FILLCELL_X2 FILLER_52_1187 ();
 FILLCELL_X4 FILLER_52_1192 ();
 FILLCELL_X2 FILLER_52_1196 ();
 FILLCELL_X8 FILLER_52_1201 ();
 FILLCELL_X16 FILLER_53_1 ();
 FILLCELL_X8 FILLER_53_20 ();
 FILLCELL_X4 FILLER_53_28 ();
 FILLCELL_X2 FILLER_53_32 ();
 FILLCELL_X2 FILLER_53_37 ();
 FILLCELL_X2 FILLER_53_42 ();
 FILLCELL_X4 FILLER_53_54 ();
 FILLCELL_X1 FILLER_53_58 ();
 FILLCELL_X1 FILLER_53_89 ();
 FILLCELL_X1 FILLER_53_113 ();
 FILLCELL_X2 FILLER_53_121 ();
 FILLCELL_X1 FILLER_53_127 ();
 FILLCELL_X4 FILLER_53_137 ();
 FILLCELL_X2 FILLER_53_141 ();
 FILLCELL_X1 FILLER_53_143 ();
 FILLCELL_X2 FILLER_53_147 ();
 FILLCELL_X2 FILLER_53_157 ();
 FILLCELL_X1 FILLER_53_159 ();
 FILLCELL_X1 FILLER_53_164 ();
 FILLCELL_X1 FILLER_53_172 ();
 FILLCELL_X2 FILLER_53_177 ();
 FILLCELL_X1 FILLER_53_179 ();
 FILLCELL_X32 FILLER_53_194 ();
 FILLCELL_X16 FILLER_53_226 ();
 FILLCELL_X8 FILLER_53_242 ();
 FILLCELL_X2 FILLER_53_250 ();
 FILLCELL_X1 FILLER_53_252 ();
 FILLCELL_X4 FILLER_53_260 ();
 FILLCELL_X2 FILLER_53_264 ();
 FILLCELL_X1 FILLER_53_301 ();
 FILLCELL_X1 FILLER_53_305 ();
 FILLCELL_X2 FILLER_53_311 ();
 FILLCELL_X1 FILLER_53_317 ();
 FILLCELL_X2 FILLER_53_321 ();
 FILLCELL_X2 FILLER_53_334 ();
 FILLCELL_X2 FILLER_53_340 ();
 FILLCELL_X1 FILLER_53_342 ();
 FILLCELL_X1 FILLER_53_361 ();
 FILLCELL_X1 FILLER_53_398 ();
 FILLCELL_X1 FILLER_53_404 ();
 FILLCELL_X4 FILLER_53_418 ();
 FILLCELL_X32 FILLER_53_428 ();
 FILLCELL_X8 FILLER_53_460 ();
 FILLCELL_X4 FILLER_53_468 ();
 FILLCELL_X1 FILLER_53_472 ();
 FILLCELL_X4 FILLER_53_485 ();
 FILLCELL_X1 FILLER_53_489 ();
 FILLCELL_X16 FILLER_53_509 ();
 FILLCELL_X4 FILLER_53_525 ();
 FILLCELL_X1 FILLER_53_529 ();
 FILLCELL_X1 FILLER_53_557 ();
 FILLCELL_X1 FILLER_53_562 ();
 FILLCELL_X1 FILLER_53_572 ();
 FILLCELL_X1 FILLER_53_634 ();
 FILLCELL_X16 FILLER_53_643 ();
 FILLCELL_X8 FILLER_53_659 ();
 FILLCELL_X2 FILLER_53_667 ();
 FILLCELL_X2 FILLER_53_672 ();
 FILLCELL_X2 FILLER_53_682 ();
 FILLCELL_X4 FILLER_53_693 ();
 FILLCELL_X2 FILLER_53_702 ();
 FILLCELL_X2 FILLER_53_720 ();
 FILLCELL_X8 FILLER_53_726 ();
 FILLCELL_X4 FILLER_53_745 ();
 FILLCELL_X1 FILLER_53_749 ();
 FILLCELL_X8 FILLER_53_754 ();
 FILLCELL_X2 FILLER_53_762 ();
 FILLCELL_X1 FILLER_53_764 ();
 FILLCELL_X1 FILLER_53_769 ();
 FILLCELL_X2 FILLER_53_774 ();
 FILLCELL_X1 FILLER_53_776 ();
 FILLCELL_X16 FILLER_53_817 ();
 FILLCELL_X1 FILLER_53_833 ();
 FILLCELL_X16 FILLER_53_860 ();
 FILLCELL_X4 FILLER_53_876 ();
 FILLCELL_X2 FILLER_53_880 ();
 FILLCELL_X1 FILLER_53_882 ();
 FILLCELL_X8 FILLER_53_896 ();
 FILLCELL_X4 FILLER_53_904 ();
 FILLCELL_X1 FILLER_53_908 ();
 FILLCELL_X8 FILLER_53_922 ();
 FILLCELL_X4 FILLER_53_930 ();
 FILLCELL_X1 FILLER_53_934 ();
 FILLCELL_X1 FILLER_53_941 ();
 FILLCELL_X1 FILLER_53_969 ();
 FILLCELL_X2 FILLER_53_976 ();
 FILLCELL_X8 FILLER_53_987 ();
 FILLCELL_X8 FILLER_53_1002 ();
 FILLCELL_X1 FILLER_53_1010 ();
 FILLCELL_X2 FILLER_53_1050 ();
 FILLCELL_X1 FILLER_53_1059 ();
 FILLCELL_X2 FILLER_53_1077 ();
 FILLCELL_X2 FILLER_53_1083 ();
 FILLCELL_X1 FILLER_53_1085 ();
 FILLCELL_X16 FILLER_53_1090 ();
 FILLCELL_X2 FILLER_53_1110 ();
 FILLCELL_X1 FILLER_53_1112 ();
 FILLCELL_X4 FILLER_53_1118 ();
 FILLCELL_X1 FILLER_53_1122 ();
 FILLCELL_X8 FILLER_53_1132 ();
 FILLCELL_X2 FILLER_53_1140 ();
 FILLCELL_X1 FILLER_53_1142 ();
 FILLCELL_X4 FILLER_53_1146 ();
 FILLCELL_X2 FILLER_53_1150 ();
 FILLCELL_X1 FILLER_53_1152 ();
 FILLCELL_X1 FILLER_53_1157 ();
 FILLCELL_X1 FILLER_53_1162 ();
 FILLCELL_X8 FILLER_53_1188 ();
 FILLCELL_X4 FILLER_53_1196 ();
 FILLCELL_X2 FILLER_53_1200 ();
 FILLCELL_X1 FILLER_53_1202 ();
 FILLCELL_X2 FILLER_53_1206 ();
 FILLCELL_X1 FILLER_53_1208 ();
 FILLCELL_X32 FILLER_54_1 ();
 FILLCELL_X4 FILLER_54_33 ();
 FILLCELL_X1 FILLER_54_37 ();
 FILLCELL_X2 FILLER_54_63 ();
 FILLCELL_X1 FILLER_54_82 ();
 FILLCELL_X1 FILLER_54_103 ();
 FILLCELL_X4 FILLER_54_115 ();
 FILLCELL_X2 FILLER_54_119 ();
 FILLCELL_X1 FILLER_54_121 ();
 FILLCELL_X2 FILLER_54_126 ();
 FILLCELL_X1 FILLER_54_128 ();
 FILLCELL_X2 FILLER_54_138 ();
 FILLCELL_X4 FILLER_54_149 ();
 FILLCELL_X2 FILLER_54_160 ();
 FILLCELL_X1 FILLER_54_162 ();
 FILLCELL_X1 FILLER_54_167 ();
 FILLCELL_X2 FILLER_54_177 ();
 FILLCELL_X1 FILLER_54_179 ();
 FILLCELL_X2 FILLER_54_184 ();
 FILLCELL_X8 FILLER_54_191 ();
 FILLCELL_X4 FILLER_54_199 ();
 FILLCELL_X4 FILLER_54_208 ();
 FILLCELL_X1 FILLER_54_212 ();
 FILLCELL_X8 FILLER_54_218 ();
 FILLCELL_X2 FILLER_54_226 ();
 FILLCELL_X1 FILLER_54_228 ();
 FILLCELL_X2 FILLER_54_246 ();
 FILLCELL_X1 FILLER_54_248 ();
 FILLCELL_X4 FILLER_54_254 ();
 FILLCELL_X4 FILLER_54_274 ();
 FILLCELL_X1 FILLER_54_308 ();
 FILLCELL_X8 FILLER_54_331 ();
 FILLCELL_X1 FILLER_54_339 ();
 FILLCELL_X16 FILLER_54_344 ();
 FILLCELL_X8 FILLER_54_360 ();
 FILLCELL_X1 FILLER_54_368 ();
 FILLCELL_X8 FILLER_54_382 ();
 FILLCELL_X2 FILLER_54_390 ();
 FILLCELL_X1 FILLER_54_392 ();
 FILLCELL_X8 FILLER_54_398 ();
 FILLCELL_X2 FILLER_54_406 ();
 FILLCELL_X2 FILLER_54_411 ();
 FILLCELL_X1 FILLER_54_413 ();
 FILLCELL_X16 FILLER_54_437 ();
 FILLCELL_X8 FILLER_54_453 ();
 FILLCELL_X4 FILLER_54_461 ();
 FILLCELL_X2 FILLER_54_465 ();
 FILLCELL_X1 FILLER_54_474 ();
 FILLCELL_X1 FILLER_54_497 ();
 FILLCELL_X8 FILLER_54_504 ();
 FILLCELL_X1 FILLER_54_537 ();
 FILLCELL_X2 FILLER_54_578 ();
 FILLCELL_X2 FILLER_54_618 ();
 FILLCELL_X1 FILLER_54_620 ();
 FILLCELL_X16 FILLER_54_635 ();
 FILLCELL_X4 FILLER_54_651 ();
 FILLCELL_X8 FILLER_54_677 ();
 FILLCELL_X1 FILLER_54_685 ();
 FILLCELL_X8 FILLER_54_689 ();
 FILLCELL_X4 FILLER_54_697 ();
 FILLCELL_X1 FILLER_54_701 ();
 FILLCELL_X4 FILLER_54_706 ();
 FILLCELL_X2 FILLER_54_710 ();
 FILLCELL_X4 FILLER_54_715 ();
 FILLCELL_X2 FILLER_54_722 ();
 FILLCELL_X1 FILLER_54_724 ();
 FILLCELL_X8 FILLER_54_739 ();
 FILLCELL_X2 FILLER_54_747 ();
 FILLCELL_X8 FILLER_54_771 ();
 FILLCELL_X2 FILLER_54_779 ();
 FILLCELL_X4 FILLER_54_800 ();
 FILLCELL_X2 FILLER_54_804 ();
 FILLCELL_X16 FILLER_54_839 ();
 FILLCELL_X2 FILLER_54_855 ();
 FILLCELL_X1 FILLER_54_857 ();
 FILLCELL_X16 FILLER_54_865 ();
 FILLCELL_X4 FILLER_54_881 ();
 FILLCELL_X2 FILLER_54_885 ();
 FILLCELL_X1 FILLER_54_904 ();
 FILLCELL_X1 FILLER_54_912 ();
 FILLCELL_X1 FILLER_54_916 ();
 FILLCELL_X8 FILLER_54_926 ();
 FILLCELL_X4 FILLER_54_934 ();
 FILLCELL_X1 FILLER_54_969 ();
 FILLCELL_X1 FILLER_54_987 ();
 FILLCELL_X2 FILLER_54_991 ();
 FILLCELL_X1 FILLER_54_995 ();
 FILLCELL_X8 FILLER_54_1005 ();
 FILLCELL_X2 FILLER_54_1013 ();
 FILLCELL_X1 FILLER_54_1015 ();
 FILLCELL_X8 FILLER_54_1019 ();
 FILLCELL_X4 FILLER_54_1027 ();
 FILLCELL_X1 FILLER_54_1031 ();
 FILLCELL_X16 FILLER_54_1034 ();
 FILLCELL_X4 FILLER_54_1050 ();
 FILLCELL_X2 FILLER_54_1054 ();
 FILLCELL_X4 FILLER_54_1060 ();
 FILLCELL_X2 FILLER_54_1064 ();
 FILLCELL_X1 FILLER_54_1078 ();
 FILLCELL_X1 FILLER_54_1083 ();
 FILLCELL_X2 FILLER_54_1107 ();
 FILLCELL_X8 FILLER_54_1121 ();
 FILLCELL_X4 FILLER_54_1129 ();
 FILLCELL_X2 FILLER_54_1133 ();
 FILLCELL_X1 FILLER_54_1135 ();
 FILLCELL_X1 FILLER_54_1147 ();
 FILLCELL_X4 FILLER_54_1164 ();
 FILLCELL_X1 FILLER_54_1168 ();
 FILLCELL_X2 FILLER_54_1181 ();
 FILLCELL_X2 FILLER_54_1191 ();
 FILLCELL_X8 FILLER_54_1196 ();
 FILLCELL_X4 FILLER_54_1204 ();
 FILLCELL_X1 FILLER_54_1208 ();
 FILLCELL_X16 FILLER_55_1 ();
 FILLCELL_X4 FILLER_55_17 ();
 FILLCELL_X16 FILLER_55_24 ();
 FILLCELL_X8 FILLER_55_40 ();
 FILLCELL_X4 FILLER_55_48 ();
 FILLCELL_X2 FILLER_55_52 ();
 FILLCELL_X4 FILLER_55_64 ();
 FILLCELL_X1 FILLER_55_68 ();
 FILLCELL_X2 FILLER_55_82 ();
 FILLCELL_X2 FILLER_55_95 ();
 FILLCELL_X1 FILLER_55_122 ();
 FILLCELL_X1 FILLER_55_134 ();
 FILLCELL_X4 FILLER_55_146 ();
 FILLCELL_X4 FILLER_55_154 ();
 FILLCELL_X2 FILLER_55_158 ();
 FILLCELL_X1 FILLER_55_160 ();
 FILLCELL_X4 FILLER_55_166 ();
 FILLCELL_X1 FILLER_55_170 ();
 FILLCELL_X16 FILLER_55_204 ();
 FILLCELL_X4 FILLER_55_220 ();
 FILLCELL_X1 FILLER_55_224 ();
 FILLCELL_X16 FILLER_55_238 ();
 FILLCELL_X2 FILLER_55_257 ();
 FILLCELL_X1 FILLER_55_297 ();
 FILLCELL_X4 FILLER_55_351 ();
 FILLCELL_X2 FILLER_55_355 ();
 FILLCELL_X1 FILLER_55_357 ();
 FILLCELL_X4 FILLER_55_368 ();
 FILLCELL_X1 FILLER_55_372 ();
 FILLCELL_X8 FILLER_55_392 ();
 FILLCELL_X4 FILLER_55_400 ();
 FILLCELL_X2 FILLER_55_404 ();
 FILLCELL_X1 FILLER_55_406 ();
 FILLCELL_X16 FILLER_55_424 ();
 FILLCELL_X8 FILLER_55_440 ();
 FILLCELL_X4 FILLER_55_448 ();
 FILLCELL_X2 FILLER_55_452 ();
 FILLCELL_X8 FILLER_55_481 ();
 FILLCELL_X2 FILLER_55_489 ();
 FILLCELL_X4 FILLER_55_501 ();
 FILLCELL_X1 FILLER_55_511 ();
 FILLCELL_X2 FILLER_55_522 ();
 FILLCELL_X1 FILLER_55_524 ();
 FILLCELL_X1 FILLER_55_549 ();
 FILLCELL_X2 FILLER_55_579 ();
 FILLCELL_X2 FILLER_55_597 ();
 FILLCELL_X1 FILLER_55_616 ();
 FILLCELL_X16 FILLER_55_625 ();
 FILLCELL_X8 FILLER_55_641 ();
 FILLCELL_X1 FILLER_55_649 ();
 FILLCELL_X8 FILLER_55_670 ();
 FILLCELL_X2 FILLER_55_678 ();
 FILLCELL_X1 FILLER_55_680 ();
 FILLCELL_X4 FILLER_55_700 ();
 FILLCELL_X1 FILLER_55_704 ();
 FILLCELL_X8 FILLER_55_719 ();
 FILLCELL_X2 FILLER_55_727 ();
 FILLCELL_X1 FILLER_55_729 ();
 FILLCELL_X8 FILLER_55_745 ();
 FILLCELL_X1 FILLER_55_766 ();
 FILLCELL_X4 FILLER_55_779 ();
 FILLCELL_X2 FILLER_55_783 ();
 FILLCELL_X1 FILLER_55_785 ();
 FILLCELL_X4 FILLER_55_814 ();
 FILLCELL_X1 FILLER_55_818 ();
 FILLCELL_X16 FILLER_55_826 ();
 FILLCELL_X8 FILLER_55_842 ();
 FILLCELL_X2 FILLER_55_850 ();
 FILLCELL_X2 FILLER_55_864 ();
 FILLCELL_X1 FILLER_55_866 ();
 FILLCELL_X1 FILLER_55_890 ();
 FILLCELL_X1 FILLER_55_898 ();
 FILLCELL_X1 FILLER_55_901 ();
 FILLCELL_X1 FILLER_55_908 ();
 FILLCELL_X1 FILLER_55_912 ();
 FILLCELL_X1 FILLER_55_916 ();
 FILLCELL_X2 FILLER_55_924 ();
 FILLCELL_X2 FILLER_55_958 ();
 FILLCELL_X1 FILLER_55_960 ();
 FILLCELL_X4 FILLER_55_970 ();
 FILLCELL_X1 FILLER_55_980 ();
 FILLCELL_X2 FILLER_55_996 ();
 FILLCELL_X1 FILLER_55_998 ();
 FILLCELL_X1 FILLER_55_1012 ();
 FILLCELL_X1 FILLER_55_1022 ();
 FILLCELL_X2 FILLER_55_1036 ();
 FILLCELL_X1 FILLER_55_1038 ();
 FILLCELL_X4 FILLER_55_1043 ();
 FILLCELL_X4 FILLER_55_1054 ();
 FILLCELL_X1 FILLER_55_1058 ();
 FILLCELL_X8 FILLER_55_1079 ();
 FILLCELL_X2 FILLER_55_1087 ();
 FILLCELL_X1 FILLER_55_1089 ();
 FILLCELL_X4 FILLER_55_1106 ();
 FILLCELL_X1 FILLER_55_1110 ();
 FILLCELL_X2 FILLER_55_1115 ();
 FILLCELL_X1 FILLER_55_1117 ();
 FILLCELL_X2 FILLER_55_1132 ();
 FILLCELL_X2 FILLER_55_1143 ();
 FILLCELL_X2 FILLER_55_1151 ();
 FILLCELL_X1 FILLER_55_1158 ();
 FILLCELL_X4 FILLER_55_1167 ();
 FILLCELL_X2 FILLER_55_1171 ();
 FILLCELL_X2 FILLER_55_1180 ();
 FILLCELL_X8 FILLER_55_1197 ();
 FILLCELL_X1 FILLER_55_1205 ();
 FILLCELL_X4 FILLER_56_1 ();
 FILLCELL_X16 FILLER_56_8 ();
 FILLCELL_X16 FILLER_56_27 ();
 FILLCELL_X4 FILLER_56_43 ();
 FILLCELL_X4 FILLER_56_67 ();
 FILLCELL_X2 FILLER_56_71 ();
 FILLCELL_X2 FILLER_56_84 ();
 FILLCELL_X2 FILLER_56_130 ();
 FILLCELL_X1 FILLER_56_136 ();
 FILLCELL_X2 FILLER_56_145 ();
 FILLCELL_X1 FILLER_56_147 ();
 FILLCELL_X4 FILLER_56_154 ();
 FILLCELL_X1 FILLER_56_158 ();
 FILLCELL_X4 FILLER_56_181 ();
 FILLCELL_X2 FILLER_56_185 ();
 FILLCELL_X16 FILLER_56_195 ();
 FILLCELL_X8 FILLER_56_211 ();
 FILLCELL_X2 FILLER_56_219 ();
 FILLCELL_X1 FILLER_56_221 ();
 FILLCELL_X16 FILLER_56_231 ();
 FILLCELL_X8 FILLER_56_247 ();
 FILLCELL_X4 FILLER_56_255 ();
 FILLCELL_X2 FILLER_56_259 ();
 FILLCELL_X2 FILLER_56_274 ();
 FILLCELL_X1 FILLER_56_276 ();
 FILLCELL_X16 FILLER_56_303 ();
 FILLCELL_X4 FILLER_56_319 ();
 FILLCELL_X1 FILLER_56_323 ();
 FILLCELL_X8 FILLER_56_335 ();
 FILLCELL_X4 FILLER_56_343 ();
 FILLCELL_X4 FILLER_56_380 ();
 FILLCELL_X2 FILLER_56_384 ();
 FILLCELL_X8 FILLER_56_390 ();
 FILLCELL_X1 FILLER_56_398 ();
 FILLCELL_X32 FILLER_56_425 ();
 FILLCELL_X2 FILLER_56_457 ();
 FILLCELL_X1 FILLER_56_467 ();
 FILLCELL_X8 FILLER_56_481 ();
 FILLCELL_X1 FILLER_56_489 ();
 FILLCELL_X2 FILLER_56_513 ();
 FILLCELL_X2 FILLER_56_525 ();
 FILLCELL_X1 FILLER_56_527 ();
 FILLCELL_X1 FILLER_56_545 ();
 FILLCELL_X2 FILLER_56_551 ();
 FILLCELL_X2 FILLER_56_599 ();
 FILLCELL_X1 FILLER_56_610 ();
 FILLCELL_X1 FILLER_56_618 ();
 FILLCELL_X2 FILLER_56_629 ();
 FILLCELL_X8 FILLER_56_632 ();
 FILLCELL_X4 FILLER_56_640 ();
 FILLCELL_X1 FILLER_56_644 ();
 FILLCELL_X2 FILLER_56_652 ();
 FILLCELL_X2 FILLER_56_658 ();
 FILLCELL_X1 FILLER_56_660 ();
 FILLCELL_X1 FILLER_56_669 ();
 FILLCELL_X2 FILLER_56_674 ();
 FILLCELL_X1 FILLER_56_676 ();
 FILLCELL_X1 FILLER_56_682 ();
 FILLCELL_X2 FILLER_56_686 ();
 FILLCELL_X1 FILLER_56_688 ();
 FILLCELL_X4 FILLER_56_704 ();
 FILLCELL_X2 FILLER_56_708 ();
 FILLCELL_X1 FILLER_56_721 ();
 FILLCELL_X2 FILLER_56_726 ();
 FILLCELL_X2 FILLER_56_732 ();
 FILLCELL_X1 FILLER_56_741 ();
 FILLCELL_X8 FILLER_56_748 ();
 FILLCELL_X4 FILLER_56_759 ();
 FILLCELL_X2 FILLER_56_763 ();
 FILLCELL_X16 FILLER_56_778 ();
 FILLCELL_X1 FILLER_56_815 ();
 FILLCELL_X16 FILLER_56_826 ();
 FILLCELL_X4 FILLER_56_842 ();
 FILLCELL_X1 FILLER_56_846 ();
 FILLCELL_X8 FILLER_56_879 ();
 FILLCELL_X16 FILLER_56_921 ();
 FILLCELL_X8 FILLER_56_937 ();
 FILLCELL_X1 FILLER_56_945 ();
 FILLCELL_X8 FILLER_56_958 ();
 FILLCELL_X1 FILLER_56_966 ();
 FILLCELL_X2 FILLER_56_979 ();
 FILLCELL_X2 FILLER_56_984 ();
 FILLCELL_X2 FILLER_56_995 ();
 FILLCELL_X1 FILLER_56_1010 ();
 FILLCELL_X4 FILLER_56_1021 ();
 FILLCELL_X1 FILLER_56_1025 ();
 FILLCELL_X32 FILLER_56_1033 ();
 FILLCELL_X4 FILLER_56_1065 ();
 FILLCELL_X2 FILLER_56_1069 ();
 FILLCELL_X2 FILLER_56_1113 ();
 FILLCELL_X2 FILLER_56_1136 ();
 FILLCELL_X4 FILLER_56_1140 ();
 FILLCELL_X2 FILLER_56_1144 ();
 FILLCELL_X1 FILLER_56_1146 ();
 FILLCELL_X16 FILLER_56_1152 ();
 FILLCELL_X16 FILLER_56_1171 ();
 FILLCELL_X4 FILLER_56_1187 ();
 FILLCELL_X2 FILLER_56_1191 ();
 FILLCELL_X1 FILLER_56_1193 ();
 FILLCELL_X4 FILLER_56_1197 ();
 FILLCELL_X2 FILLER_56_1201 ();
 FILLCELL_X1 FILLER_56_1203 ();
 FILLCELL_X2 FILLER_56_1207 ();
 FILLCELL_X2 FILLER_57_1 ();
 FILLCELL_X1 FILLER_57_3 ();
 FILLCELL_X16 FILLER_57_7 ();
 FILLCELL_X32 FILLER_57_26 ();
 FILLCELL_X8 FILLER_57_58 ();
 FILLCELL_X4 FILLER_57_75 ();
 FILLCELL_X2 FILLER_57_79 ();
 FILLCELL_X1 FILLER_57_100 ();
 FILLCELL_X4 FILLER_57_135 ();
 FILLCELL_X2 FILLER_57_139 ();
 FILLCELL_X1 FILLER_57_141 ();
 FILLCELL_X4 FILLER_57_156 ();
 FILLCELL_X1 FILLER_57_160 ();
 FILLCELL_X1 FILLER_57_165 ();
 FILLCELL_X1 FILLER_57_177 ();
 FILLCELL_X4 FILLER_57_182 ();
 FILLCELL_X2 FILLER_57_186 ();
 FILLCELL_X8 FILLER_57_195 ();
 FILLCELL_X1 FILLER_57_203 ();
 FILLCELL_X4 FILLER_57_221 ();
 FILLCELL_X2 FILLER_57_225 ();
 FILLCELL_X1 FILLER_57_227 ();
 FILLCELL_X4 FILLER_57_245 ();
 FILLCELL_X1 FILLER_57_249 ();
 FILLCELL_X1 FILLER_57_272 ();
 FILLCELL_X4 FILLER_57_309 ();
 FILLCELL_X4 FILLER_57_326 ();
 FILLCELL_X1 FILLER_57_359 ();
 FILLCELL_X1 FILLER_57_365 ();
 FILLCELL_X8 FILLER_57_390 ();
 FILLCELL_X2 FILLER_57_398 ();
 FILLCELL_X2 FILLER_57_415 ();
 FILLCELL_X16 FILLER_57_425 ();
 FILLCELL_X8 FILLER_57_441 ();
 FILLCELL_X4 FILLER_57_449 ();
 FILLCELL_X2 FILLER_57_453 ();
 FILLCELL_X4 FILLER_57_525 ();
 FILLCELL_X1 FILLER_57_529 ();
 FILLCELL_X16 FILLER_57_537 ();
 FILLCELL_X4 FILLER_57_553 ();
 FILLCELL_X1 FILLER_57_557 ();
 FILLCELL_X2 FILLER_57_599 ();
 FILLCELL_X8 FILLER_57_608 ();
 FILLCELL_X2 FILLER_57_616 ();
 FILLCELL_X1 FILLER_57_624 ();
 FILLCELL_X16 FILLER_57_635 ();
 FILLCELL_X2 FILLER_57_651 ();
 FILLCELL_X1 FILLER_57_653 ();
 FILLCELL_X1 FILLER_57_658 ();
 FILLCELL_X4 FILLER_57_663 ();
 FILLCELL_X1 FILLER_57_667 ();
 FILLCELL_X8 FILLER_57_672 ();
 FILLCELL_X2 FILLER_57_680 ();
 FILLCELL_X16 FILLER_57_685 ();
 FILLCELL_X2 FILLER_57_701 ();
 FILLCELL_X1 FILLER_57_703 ();
 FILLCELL_X8 FILLER_57_724 ();
 FILLCELL_X4 FILLER_57_732 ();
 FILLCELL_X1 FILLER_57_736 ();
 FILLCELL_X8 FILLER_57_741 ();
 FILLCELL_X2 FILLER_57_749 ();
 FILLCELL_X1 FILLER_57_751 ();
 FILLCELL_X4 FILLER_57_759 ();
 FILLCELL_X2 FILLER_57_763 ();
 FILLCELL_X1 FILLER_57_765 ();
 FILLCELL_X2 FILLER_57_770 ();
 FILLCELL_X1 FILLER_57_772 ();
 FILLCELL_X2 FILLER_57_775 ();
 FILLCELL_X1 FILLER_57_777 ();
 FILLCELL_X2 FILLER_57_781 ();
 FILLCELL_X1 FILLER_57_783 ();
 FILLCELL_X1 FILLER_57_788 ();
 FILLCELL_X1 FILLER_57_796 ();
 FILLCELL_X2 FILLER_57_801 ();
 FILLCELL_X4 FILLER_57_807 ();
 FILLCELL_X2 FILLER_57_811 ();
 FILLCELL_X32 FILLER_57_817 ();
 FILLCELL_X4 FILLER_57_849 ();
 FILLCELL_X2 FILLER_57_853 ();
 FILLCELL_X4 FILLER_57_879 ();
 FILLCELL_X2 FILLER_57_883 ();
 FILLCELL_X1 FILLER_57_885 ();
 FILLCELL_X1 FILLER_57_892 ();
 FILLCELL_X1 FILLER_57_896 ();
 FILLCELL_X4 FILLER_57_904 ();
 FILLCELL_X1 FILLER_57_908 ();
 FILLCELL_X2 FILLER_57_918 ();
 FILLCELL_X1 FILLER_57_935 ();
 FILLCELL_X4 FILLER_57_946 ();
 FILLCELL_X1 FILLER_57_950 ();
 FILLCELL_X4 FILLER_57_957 ();
 FILLCELL_X2 FILLER_57_961 ();
 FILLCELL_X4 FILLER_57_983 ();
 FILLCELL_X2 FILLER_57_987 ();
 FILLCELL_X1 FILLER_57_989 ();
 FILLCELL_X8 FILLER_57_1009 ();
 FILLCELL_X4 FILLER_57_1017 ();
 FILLCELL_X2 FILLER_57_1021 ();
 FILLCELL_X1 FILLER_57_1023 ();
 FILLCELL_X32 FILLER_57_1043 ();
 FILLCELL_X32 FILLER_57_1075 ();
 FILLCELL_X16 FILLER_57_1107 ();
 FILLCELL_X8 FILLER_57_1123 ();
 FILLCELL_X4 FILLER_57_1131 ();
 FILLCELL_X1 FILLER_57_1135 ();
 FILLCELL_X32 FILLER_57_1140 ();
 FILLCELL_X4 FILLER_57_1172 ();
 FILLCELL_X2 FILLER_57_1176 ();
 FILLCELL_X1 FILLER_57_1178 ();
 FILLCELL_X16 FILLER_57_1182 ();
 FILLCELL_X4 FILLER_57_1201 ();
 FILLCELL_X1 FILLER_57_1205 ();
 FILLCELL_X16 FILLER_58_1 ();
 FILLCELL_X4 FILLER_58_17 ();
 FILLCELL_X2 FILLER_58_21 ();
 FILLCELL_X1 FILLER_58_23 ();
 FILLCELL_X32 FILLER_58_27 ();
 FILLCELL_X4 FILLER_58_59 ();
 FILLCELL_X2 FILLER_58_63 ();
 FILLCELL_X8 FILLER_58_78 ();
 FILLCELL_X1 FILLER_58_86 ();
 FILLCELL_X2 FILLER_58_89 ();
 FILLCELL_X1 FILLER_58_105 ();
 FILLCELL_X2 FILLER_58_124 ();
 FILLCELL_X1 FILLER_58_126 ();
 FILLCELL_X8 FILLER_58_134 ();
 FILLCELL_X4 FILLER_58_142 ();
 FILLCELL_X1 FILLER_58_146 ();
 FILLCELL_X2 FILLER_58_160 ();
 FILLCELL_X2 FILLER_58_169 ();
 FILLCELL_X2 FILLER_58_182 ();
 FILLCELL_X4 FILLER_58_196 ();
 FILLCELL_X2 FILLER_58_207 ();
 FILLCELL_X2 FILLER_58_214 ();
 FILLCELL_X1 FILLER_58_219 ();
 FILLCELL_X8 FILLER_58_238 ();
 FILLCELL_X4 FILLER_58_246 ();
 FILLCELL_X2 FILLER_58_250 ();
 FILLCELL_X4 FILLER_58_316 ();
 FILLCELL_X2 FILLER_58_320 ();
 FILLCELL_X1 FILLER_58_326 ();
 FILLCELL_X4 FILLER_58_334 ();
 FILLCELL_X1 FILLER_58_338 ();
 FILLCELL_X1 FILLER_58_350 ();
 FILLCELL_X4 FILLER_58_360 ();
 FILLCELL_X2 FILLER_58_364 ();
 FILLCELL_X4 FILLER_58_370 ();
 FILLCELL_X2 FILLER_58_385 ();
 FILLCELL_X8 FILLER_58_402 ();
 FILLCELL_X1 FILLER_58_410 ();
 FILLCELL_X2 FILLER_58_423 ();
 FILLCELL_X32 FILLER_58_434 ();
 FILLCELL_X4 FILLER_58_472 ();
 FILLCELL_X2 FILLER_58_489 ();
 FILLCELL_X1 FILLER_58_491 ();
 FILLCELL_X2 FILLER_58_499 ();
 FILLCELL_X4 FILLER_58_516 ();
 FILLCELL_X1 FILLER_58_520 ();
 FILLCELL_X1 FILLER_58_527 ();
 FILLCELL_X16 FILLER_58_542 ();
 FILLCELL_X1 FILLER_58_558 ();
 FILLCELL_X1 FILLER_58_569 ();
 FILLCELL_X4 FILLER_58_591 ();
 FILLCELL_X2 FILLER_58_595 ();
 FILLCELL_X16 FILLER_58_610 ();
 FILLCELL_X4 FILLER_58_626 ();
 FILLCELL_X1 FILLER_58_630 ();
 FILLCELL_X16 FILLER_58_632 ();
 FILLCELL_X8 FILLER_58_648 ();
 FILLCELL_X4 FILLER_58_656 ();
 FILLCELL_X1 FILLER_58_660 ();
 FILLCELL_X2 FILLER_58_665 ();
 FILLCELL_X1 FILLER_58_667 ();
 FILLCELL_X2 FILLER_58_672 ();
 FILLCELL_X1 FILLER_58_674 ();
 FILLCELL_X4 FILLER_58_693 ();
 FILLCELL_X8 FILLER_58_700 ();
 FILLCELL_X4 FILLER_58_708 ();
 FILLCELL_X2 FILLER_58_712 ();
 FILLCELL_X1 FILLER_58_714 ();
 FILLCELL_X4 FILLER_58_718 ();
 FILLCELL_X8 FILLER_58_727 ();
 FILLCELL_X2 FILLER_58_745 ();
 FILLCELL_X1 FILLER_58_747 ();
 FILLCELL_X2 FILLER_58_755 ();
 FILLCELL_X8 FILLER_58_760 ();
 FILLCELL_X4 FILLER_58_773 ();
 FILLCELL_X2 FILLER_58_777 ();
 FILLCELL_X1 FILLER_58_779 ();
 FILLCELL_X1 FILLER_58_800 ();
 FILLCELL_X4 FILLER_58_809 ();
 FILLCELL_X2 FILLER_58_813 ();
 FILLCELL_X1 FILLER_58_815 ();
 FILLCELL_X16 FILLER_58_826 ();
 FILLCELL_X8 FILLER_58_842 ();
 FILLCELL_X4 FILLER_58_850 ();
 FILLCELL_X2 FILLER_58_854 ();
 FILLCELL_X1 FILLER_58_856 ();
 FILLCELL_X1 FILLER_58_863 ();
 FILLCELL_X8 FILLER_58_874 ();
 FILLCELL_X2 FILLER_58_882 ();
 FILLCELL_X1 FILLER_58_884 ();
 FILLCELL_X1 FILLER_58_894 ();
 FILLCELL_X2 FILLER_58_912 ();
 FILLCELL_X1 FILLER_58_918 ();
 FILLCELL_X2 FILLER_58_928 ();
 FILLCELL_X8 FILLER_58_936 ();
 FILLCELL_X4 FILLER_58_944 ();
 FILLCELL_X2 FILLER_58_948 ();
 FILLCELL_X1 FILLER_58_950 ();
 FILLCELL_X1 FILLER_58_969 ();
 FILLCELL_X2 FILLER_58_976 ();
 FILLCELL_X4 FILLER_58_988 ();
 FILLCELL_X2 FILLER_58_1025 ();
 FILLCELL_X16 FILLER_58_1033 ();
 FILLCELL_X4 FILLER_58_1049 ();
 FILLCELL_X2 FILLER_58_1053 ();
 FILLCELL_X16 FILLER_58_1072 ();
 FILLCELL_X4 FILLER_58_1088 ();
 FILLCELL_X1 FILLER_58_1092 ();
 FILLCELL_X1 FILLER_58_1110 ();
 FILLCELL_X8 FILLER_58_1133 ();
 FILLCELL_X32 FILLER_58_1158 ();
 FILLCELL_X4 FILLER_58_1190 ();
 FILLCELL_X8 FILLER_58_1197 ();
 FILLCELL_X4 FILLER_58_1205 ();
 FILLCELL_X16 FILLER_59_1 ();
 FILLCELL_X8 FILLER_59_17 ();
 FILLCELL_X4 FILLER_59_25 ();
 FILLCELL_X32 FILLER_59_32 ();
 FILLCELL_X2 FILLER_59_64 ();
 FILLCELL_X1 FILLER_59_66 ();
 FILLCELL_X4 FILLER_59_80 ();
 FILLCELL_X2 FILLER_59_84 ();
 FILLCELL_X1 FILLER_59_86 ();
 FILLCELL_X4 FILLER_59_101 ();
 FILLCELL_X4 FILLER_59_112 ();
 FILLCELL_X1 FILLER_59_116 ();
 FILLCELL_X2 FILLER_59_135 ();
 FILLCELL_X8 FILLER_59_151 ();
 FILLCELL_X1 FILLER_59_159 ();
 FILLCELL_X1 FILLER_59_167 ();
 FILLCELL_X1 FILLER_59_178 ();
 FILLCELL_X16 FILLER_59_191 ();
 FILLCELL_X8 FILLER_59_216 ();
 FILLCELL_X2 FILLER_59_224 ();
 FILLCELL_X2 FILLER_59_229 ();
 FILLCELL_X8 FILLER_59_240 ();
 FILLCELL_X1 FILLER_59_275 ();
 FILLCELL_X2 FILLER_59_280 ();
 FILLCELL_X1 FILLER_59_282 ();
 FILLCELL_X1 FILLER_59_297 ();
 FILLCELL_X4 FILLER_59_323 ();
 FILLCELL_X1 FILLER_59_327 ();
 FILLCELL_X16 FILLER_59_332 ();
 FILLCELL_X4 FILLER_59_348 ();
 FILLCELL_X1 FILLER_59_352 ();
 FILLCELL_X2 FILLER_59_357 ();
 FILLCELL_X4 FILLER_59_374 ();
 FILLCELL_X1 FILLER_59_378 ();
 FILLCELL_X8 FILLER_59_390 ();
 FILLCELL_X8 FILLER_59_443 ();
 FILLCELL_X4 FILLER_59_451 ();
 FILLCELL_X1 FILLER_59_455 ();
 FILLCELL_X4 FILLER_59_473 ();
 FILLCELL_X2 FILLER_59_477 ();
 FILLCELL_X1 FILLER_59_479 ();
 FILLCELL_X2 FILLER_59_511 ();
 FILLCELL_X2 FILLER_59_522 ();
 FILLCELL_X1 FILLER_59_524 ();
 FILLCELL_X8 FILLER_59_529 ();
 FILLCELL_X2 FILLER_59_537 ();
 FILLCELL_X1 FILLER_59_539 ();
 FILLCELL_X1 FILLER_59_542 ();
 FILLCELL_X2 FILLER_59_557 ();
 FILLCELL_X4 FILLER_59_565 ();
 FILLCELL_X1 FILLER_59_569 ();
 FILLCELL_X4 FILLER_59_582 ();
 FILLCELL_X2 FILLER_59_595 ();
 FILLCELL_X1 FILLER_59_597 ();
 FILLCELL_X16 FILLER_59_604 ();
 FILLCELL_X8 FILLER_59_620 ();
 FILLCELL_X4 FILLER_59_628 ();
 FILLCELL_X16 FILLER_59_636 ();
 FILLCELL_X16 FILLER_59_668 ();
 FILLCELL_X4 FILLER_59_684 ();
 FILLCELL_X2 FILLER_59_688 ();
 FILLCELL_X1 FILLER_59_690 ();
 FILLCELL_X16 FILLER_59_695 ();
 FILLCELL_X8 FILLER_59_711 ();
 FILLCELL_X4 FILLER_59_719 ();
 FILLCELL_X16 FILLER_59_732 ();
 FILLCELL_X8 FILLER_59_748 ();
 FILLCELL_X4 FILLER_59_756 ();
 FILLCELL_X4 FILLER_59_762 ();
 FILLCELL_X2 FILLER_59_766 ();
 FILLCELL_X8 FILLER_59_774 ();
 FILLCELL_X8 FILLER_59_806 ();
 FILLCELL_X1 FILLER_59_814 ();
 FILLCELL_X32 FILLER_59_819 ();
 FILLCELL_X1 FILLER_59_851 ();
 FILLCELL_X1 FILLER_59_855 ();
 FILLCELL_X1 FILLER_59_863 ();
 FILLCELL_X2 FILLER_59_873 ();
 FILLCELL_X1 FILLER_59_875 ();
 FILLCELL_X2 FILLER_59_897 ();
 FILLCELL_X1 FILLER_59_932 ();
 FILLCELL_X2 FILLER_59_951 ();
 FILLCELL_X4 FILLER_59_965 ();
 FILLCELL_X1 FILLER_59_979 ();
 FILLCELL_X1 FILLER_59_986 ();
 FILLCELL_X4 FILLER_59_1011 ();
 FILLCELL_X1 FILLER_59_1015 ();
 FILLCELL_X4 FILLER_59_1028 ();
 FILLCELL_X2 FILLER_59_1032 ();
 FILLCELL_X32 FILLER_59_1051 ();
 FILLCELL_X2 FILLER_59_1083 ();
 FILLCELL_X8 FILLER_59_1091 ();
 FILLCELL_X4 FILLER_59_1099 ();
 FILLCELL_X2 FILLER_59_1103 ();
 FILLCELL_X1 FILLER_59_1105 ();
 FILLCELL_X16 FILLER_59_1149 ();
 FILLCELL_X8 FILLER_59_1165 ();
 FILLCELL_X4 FILLER_59_1173 ();
 FILLCELL_X1 FILLER_59_1177 ();
 FILLCELL_X8 FILLER_59_1198 ();
 FILLCELL_X2 FILLER_59_1206 ();
 FILLCELL_X1 FILLER_59_1208 ();
 FILLCELL_X32 FILLER_60_1 ();
 FILLCELL_X32 FILLER_60_33 ();
 FILLCELL_X2 FILLER_60_65 ();
 FILLCELL_X1 FILLER_60_67 ();
 FILLCELL_X4 FILLER_60_77 ();
 FILLCELL_X1 FILLER_60_81 ();
 FILLCELL_X2 FILLER_60_98 ();
 FILLCELL_X1 FILLER_60_100 ();
 FILLCELL_X4 FILLER_60_108 ();
 FILLCELL_X1 FILLER_60_119 ();
 FILLCELL_X1 FILLER_60_129 ();
 FILLCELL_X1 FILLER_60_147 ();
 FILLCELL_X4 FILLER_60_175 ();
 FILLCELL_X1 FILLER_60_188 ();
 FILLCELL_X1 FILLER_60_195 ();
 FILLCELL_X4 FILLER_60_212 ();
 FILLCELL_X4 FILLER_60_237 ();
 FILLCELL_X2 FILLER_60_241 ();
 FILLCELL_X8 FILLER_60_302 ();
 FILLCELL_X2 FILLER_60_310 ();
 FILLCELL_X1 FILLER_60_312 ();
 FILLCELL_X2 FILLER_60_331 ();
 FILLCELL_X1 FILLER_60_333 ();
 FILLCELL_X8 FILLER_60_338 ();
 FILLCELL_X4 FILLER_60_351 ();
 FILLCELL_X2 FILLER_60_365 ();
 FILLCELL_X1 FILLER_60_367 ();
 FILLCELL_X1 FILLER_60_376 ();
 FILLCELL_X2 FILLER_60_385 ();
 FILLCELL_X2 FILLER_60_393 ();
 FILLCELL_X1 FILLER_60_395 ();
 FILLCELL_X1 FILLER_60_419 ();
 FILLCELL_X4 FILLER_60_428 ();
 FILLCELL_X2 FILLER_60_432 ();
 FILLCELL_X16 FILLER_60_451 ();
 FILLCELL_X1 FILLER_60_467 ();
 FILLCELL_X1 FILLER_60_492 ();
 FILLCELL_X2 FILLER_60_507 ();
 FILLCELL_X1 FILLER_60_509 ();
 FILLCELL_X1 FILLER_60_537 ();
 FILLCELL_X1 FILLER_60_556 ();
 FILLCELL_X2 FILLER_60_573 ();
 FILLCELL_X1 FILLER_60_575 ();
 FILLCELL_X2 FILLER_60_585 ();
 FILLCELL_X1 FILLER_60_587 ();
 FILLCELL_X2 FILLER_60_597 ();
 FILLCELL_X8 FILLER_60_609 ();
 FILLCELL_X4 FILLER_60_626 ();
 FILLCELL_X1 FILLER_60_630 ();
 FILLCELL_X16 FILLER_60_632 ();
 FILLCELL_X1 FILLER_60_648 ();
 FILLCELL_X1 FILLER_60_656 ();
 FILLCELL_X2 FILLER_60_665 ();
 FILLCELL_X4 FILLER_60_693 ();
 FILLCELL_X2 FILLER_60_710 ();
 FILLCELL_X1 FILLER_60_719 ();
 FILLCELL_X8 FILLER_60_729 ();
 FILLCELL_X1 FILLER_60_737 ();
 FILLCELL_X4 FILLER_60_742 ();
 FILLCELL_X2 FILLER_60_746 ();
 FILLCELL_X1 FILLER_60_748 ();
 FILLCELL_X4 FILLER_60_752 ();
 FILLCELL_X2 FILLER_60_756 ();
 FILLCELL_X1 FILLER_60_758 ();
 FILLCELL_X8 FILLER_60_773 ();
 FILLCELL_X1 FILLER_60_781 ();
 FILLCELL_X4 FILLER_60_786 ();
 FILLCELL_X4 FILLER_60_802 ();
 FILLCELL_X2 FILLER_60_819 ();
 FILLCELL_X8 FILLER_60_826 ();
 FILLCELL_X4 FILLER_60_853 ();
 FILLCELL_X1 FILLER_60_857 ();
 FILLCELL_X1 FILLER_60_861 ();
 FILLCELL_X2 FILLER_60_883 ();
 FILLCELL_X1 FILLER_60_885 ();
 FILLCELL_X1 FILLER_60_906 ();
 FILLCELL_X2 FILLER_60_939 ();
 FILLCELL_X1 FILLER_60_941 ();
 FILLCELL_X2 FILLER_60_962 ();
 FILLCELL_X8 FILLER_60_989 ();
 FILLCELL_X4 FILLER_60_997 ();
 FILLCELL_X1 FILLER_60_1001 ();
 FILLCELL_X16 FILLER_60_1011 ();
 FILLCELL_X8 FILLER_60_1027 ();
 FILLCELL_X2 FILLER_60_1035 ();
 FILLCELL_X1 FILLER_60_1037 ();
 FILLCELL_X4 FILLER_60_1068 ();
 FILLCELL_X8 FILLER_60_1082 ();
 FILLCELL_X1 FILLER_60_1090 ();
 FILLCELL_X2 FILLER_60_1112 ();
 FILLCELL_X8 FILLER_60_1124 ();
 FILLCELL_X4 FILLER_60_1132 ();
 FILLCELL_X2 FILLER_60_1136 ();
 FILLCELL_X8 FILLER_60_1153 ();
 FILLCELL_X2 FILLER_60_1161 ();
 FILLCELL_X1 FILLER_60_1163 ();
 FILLCELL_X2 FILLER_60_1168 ();
 FILLCELL_X1 FILLER_60_1170 ();
 FILLCELL_X2 FILLER_60_1188 ();
 FILLCELL_X1 FILLER_60_1190 ();
 FILLCELL_X4 FILLER_60_1194 ();
 FILLCELL_X2 FILLER_60_1198 ();
 FILLCELL_X1 FILLER_60_1200 ();
 FILLCELL_X4 FILLER_60_1204 ();
 FILLCELL_X1 FILLER_60_1208 ();
 FILLCELL_X16 FILLER_61_1 ();
 FILLCELL_X4 FILLER_61_17 ();
 FILLCELL_X2 FILLER_61_21 ();
 FILLCELL_X1 FILLER_61_23 ();
 FILLCELL_X32 FILLER_61_27 ();
 FILLCELL_X16 FILLER_61_59 ();
 FILLCELL_X4 FILLER_61_75 ();
 FILLCELL_X4 FILLER_61_92 ();
 FILLCELL_X2 FILLER_61_96 ();
 FILLCELL_X2 FILLER_61_105 ();
 FILLCELL_X1 FILLER_61_107 ();
 FILLCELL_X2 FILLER_61_133 ();
 FILLCELL_X2 FILLER_61_149 ();
 FILLCELL_X4 FILLER_61_158 ();
 FILLCELL_X1 FILLER_61_162 ();
 FILLCELL_X1 FILLER_61_171 ();
 FILLCELL_X16 FILLER_61_191 ();
 FILLCELL_X8 FILLER_61_207 ();
 FILLCELL_X16 FILLER_61_232 ();
 FILLCELL_X4 FILLER_61_248 ();
 FILLCELL_X2 FILLER_61_278 ();
 FILLCELL_X1 FILLER_61_284 ();
 FILLCELL_X2 FILLER_61_292 ();
 FILLCELL_X2 FILLER_61_298 ();
 FILLCELL_X2 FILLER_61_307 ();
 FILLCELL_X1 FILLER_61_309 ();
 FILLCELL_X2 FILLER_61_314 ();
 FILLCELL_X1 FILLER_61_316 ();
 FILLCELL_X2 FILLER_61_321 ();
 FILLCELL_X1 FILLER_61_333 ();
 FILLCELL_X2 FILLER_61_345 ();
 FILLCELL_X1 FILLER_61_361 ();
 FILLCELL_X2 FILLER_61_367 ();
 FILLCELL_X1 FILLER_61_369 ();
 FILLCELL_X1 FILLER_61_379 ();
 FILLCELL_X4 FILLER_61_399 ();
 FILLCELL_X1 FILLER_61_403 ();
 FILLCELL_X1 FILLER_61_408 ();
 FILLCELL_X32 FILLER_61_424 ();
 FILLCELL_X16 FILLER_61_456 ();
 FILLCELL_X8 FILLER_61_472 ();
 FILLCELL_X1 FILLER_61_480 ();
 FILLCELL_X1 FILLER_61_484 ();
 FILLCELL_X8 FILLER_61_519 ();
 FILLCELL_X1 FILLER_61_527 ();
 FILLCELL_X4 FILLER_61_547 ();
 FILLCELL_X2 FILLER_61_554 ();
 FILLCELL_X1 FILLER_61_556 ();
 FILLCELL_X2 FILLER_61_560 ();
 FILLCELL_X1 FILLER_61_562 ();
 FILLCELL_X2 FILLER_61_576 ();
 FILLCELL_X8 FILLER_61_607 ();
 FILLCELL_X4 FILLER_61_615 ();
 FILLCELL_X1 FILLER_61_619 ();
 FILLCELL_X8 FILLER_61_637 ();
 FILLCELL_X4 FILLER_61_665 ();
 FILLCELL_X1 FILLER_61_669 ();
 FILLCELL_X4 FILLER_61_677 ();
 FILLCELL_X1 FILLER_61_681 ();
 FILLCELL_X4 FILLER_61_688 ();
 FILLCELL_X2 FILLER_61_692 ();
 FILLCELL_X1 FILLER_61_694 ();
 FILLCELL_X8 FILLER_61_700 ();
 FILLCELL_X4 FILLER_61_708 ();
 FILLCELL_X2 FILLER_61_719 ();
 FILLCELL_X1 FILLER_61_721 ();
 FILLCELL_X2 FILLER_61_729 ();
 FILLCELL_X1 FILLER_61_731 ();
 FILLCELL_X16 FILLER_61_741 ();
 FILLCELL_X4 FILLER_61_757 ();
 FILLCELL_X2 FILLER_61_767 ();
 FILLCELL_X4 FILLER_61_776 ();
 FILLCELL_X1 FILLER_61_780 ();
 FILLCELL_X1 FILLER_61_792 ();
 FILLCELL_X2 FILLER_61_810 ();
 FILLCELL_X1 FILLER_61_812 ();
 FILLCELL_X2 FILLER_61_881 ();
 FILLCELL_X1 FILLER_61_883 ();
 FILLCELL_X2 FILLER_61_896 ();
 FILLCELL_X1 FILLER_61_898 ();
 FILLCELL_X2 FILLER_61_929 ();
 FILLCELL_X1 FILLER_61_931 ();
 FILLCELL_X2 FILLER_61_950 ();
 FILLCELL_X2 FILLER_61_976 ();
 FILLCELL_X1 FILLER_61_981 ();
 FILLCELL_X1 FILLER_61_992 ();
 FILLCELL_X16 FILLER_61_996 ();
 FILLCELL_X8 FILLER_61_1012 ();
 FILLCELL_X4 FILLER_61_1020 ();
 FILLCELL_X2 FILLER_61_1024 ();
 FILLCELL_X1 FILLER_61_1026 ();
 FILLCELL_X2 FILLER_61_1066 ();
 FILLCELL_X1 FILLER_61_1077 ();
 FILLCELL_X8 FILLER_61_1093 ();
 FILLCELL_X1 FILLER_61_1101 ();
 FILLCELL_X2 FILLER_61_1112 ();
 FILLCELL_X1 FILLER_61_1154 ();
 FILLCELL_X8 FILLER_61_1197 ();
 FILLCELL_X4 FILLER_61_1205 ();
 FILLCELL_X32 FILLER_62_1 ();
 FILLCELL_X32 FILLER_62_33 ();
 FILLCELL_X32 FILLER_62_65 ();
 FILLCELL_X2 FILLER_62_110 ();
 FILLCELL_X1 FILLER_62_125 ();
 FILLCELL_X1 FILLER_62_143 ();
 FILLCELL_X2 FILLER_62_151 ();
 FILLCELL_X2 FILLER_62_165 ();
 FILLCELL_X1 FILLER_62_177 ();
 FILLCELL_X8 FILLER_62_191 ();
 FILLCELL_X4 FILLER_62_199 ();
 FILLCELL_X2 FILLER_62_203 ();
 FILLCELL_X4 FILLER_62_251 ();
 FILLCELL_X1 FILLER_62_289 ();
 FILLCELL_X2 FILLER_62_307 ();
 FILLCELL_X1 FILLER_62_313 ();
 FILLCELL_X16 FILLER_62_323 ();
 FILLCELL_X4 FILLER_62_339 ();
 FILLCELL_X4 FILLER_62_368 ();
 FILLCELL_X1 FILLER_62_372 ();
 FILLCELL_X8 FILLER_62_376 ();
 FILLCELL_X4 FILLER_62_384 ();
 FILLCELL_X4 FILLER_62_399 ();
 FILLCELL_X2 FILLER_62_403 ();
 FILLCELL_X1 FILLER_62_405 ();
 FILLCELL_X1 FILLER_62_410 ();
 FILLCELL_X2 FILLER_62_416 ();
 FILLCELL_X2 FILLER_62_422 ();
 FILLCELL_X1 FILLER_62_424 ();
 FILLCELL_X2 FILLER_62_438 ();
 FILLCELL_X1 FILLER_62_440 ();
 FILLCELL_X8 FILLER_62_450 ();
 FILLCELL_X1 FILLER_62_458 ();
 FILLCELL_X4 FILLER_62_498 ();
 FILLCELL_X1 FILLER_62_502 ();
 FILLCELL_X4 FILLER_62_564 ();
 FILLCELL_X2 FILLER_62_568 ();
 FILLCELL_X16 FILLER_62_604 ();
 FILLCELL_X8 FILLER_62_620 ();
 FILLCELL_X2 FILLER_62_628 ();
 FILLCELL_X1 FILLER_62_630 ();
 FILLCELL_X8 FILLER_62_632 ();
 FILLCELL_X4 FILLER_62_640 ();
 FILLCELL_X2 FILLER_62_644 ();
 FILLCELL_X16 FILLER_62_650 ();
 FILLCELL_X4 FILLER_62_671 ();
 FILLCELL_X16 FILLER_62_686 ();
 FILLCELL_X8 FILLER_62_702 ();
 FILLCELL_X4 FILLER_62_710 ();
 FILLCELL_X1 FILLER_62_730 ();
 FILLCELL_X1 FILLER_62_742 ();
 FILLCELL_X8 FILLER_62_749 ();
 FILLCELL_X2 FILLER_62_757 ();
 FILLCELL_X1 FILLER_62_759 ();
 FILLCELL_X2 FILLER_62_763 ();
 FILLCELL_X4 FILLER_62_776 ();
 FILLCELL_X2 FILLER_62_780 ();
 FILLCELL_X1 FILLER_62_782 ();
 FILLCELL_X2 FILLER_62_793 ();
 FILLCELL_X1 FILLER_62_801 ();
 FILLCELL_X1 FILLER_62_812 ();
 FILLCELL_X1 FILLER_62_817 ();
 FILLCELL_X4 FILLER_62_828 ();
 FILLCELL_X16 FILLER_62_841 ();
 FILLCELL_X8 FILLER_62_857 ();
 FILLCELL_X2 FILLER_62_865 ();
 FILLCELL_X1 FILLER_62_867 ();
 FILLCELL_X2 FILLER_62_895 ();
 FILLCELL_X2 FILLER_62_910 ();
 FILLCELL_X1 FILLER_62_912 ();
 FILLCELL_X8 FILLER_62_923 ();
 FILLCELL_X4 FILLER_62_931 ();
 FILLCELL_X2 FILLER_62_935 ();
 FILLCELL_X4 FILLER_62_947 ();
 FILLCELL_X2 FILLER_62_975 ();
 FILLCELL_X1 FILLER_62_977 ();
 FILLCELL_X1 FILLER_62_990 ();
 FILLCELL_X2 FILLER_62_1000 ();
 FILLCELL_X1 FILLER_62_1006 ();
 FILLCELL_X4 FILLER_62_1014 ();
 FILLCELL_X2 FILLER_62_1018 ();
 FILLCELL_X1 FILLER_62_1020 ();
 FILLCELL_X4 FILLER_62_1028 ();
 FILLCELL_X1 FILLER_62_1032 ();
 FILLCELL_X1 FILLER_62_1053 ();
 FILLCELL_X1 FILLER_62_1104 ();
 FILLCELL_X1 FILLER_62_1140 ();
 FILLCELL_X2 FILLER_62_1145 ();
 FILLCELL_X1 FILLER_62_1147 ();
 FILLCELL_X8 FILLER_62_1178 ();
 FILLCELL_X4 FILLER_62_1186 ();
 FILLCELL_X2 FILLER_62_1190 ();
 FILLCELL_X1 FILLER_62_1192 ();
 FILLCELL_X4 FILLER_62_1200 ();
 FILLCELL_X2 FILLER_62_1204 ();
 FILLCELL_X32 FILLER_63_1 ();
 FILLCELL_X8 FILLER_63_33 ();
 FILLCELL_X32 FILLER_63_49 ();
 FILLCELL_X16 FILLER_63_81 ();
 FILLCELL_X8 FILLER_63_97 ();
 FILLCELL_X4 FILLER_63_105 ();
 FILLCELL_X2 FILLER_63_109 ();
 FILLCELL_X16 FILLER_63_136 ();
 FILLCELL_X8 FILLER_63_152 ();
 FILLCELL_X4 FILLER_63_160 ();
 FILLCELL_X1 FILLER_63_164 ();
 FILLCELL_X4 FILLER_63_178 ();
 FILLCELL_X2 FILLER_63_182 ();
 FILLCELL_X1 FILLER_63_184 ();
 FILLCELL_X32 FILLER_63_188 ();
 FILLCELL_X1 FILLER_63_220 ();
 FILLCELL_X8 FILLER_63_260 ();
 FILLCELL_X2 FILLER_63_268 ();
 FILLCELL_X1 FILLER_63_270 ();
 FILLCELL_X4 FILLER_63_274 ();
 FILLCELL_X2 FILLER_63_278 ();
 FILLCELL_X1 FILLER_63_280 ();
 FILLCELL_X4 FILLER_63_307 ();
 FILLCELL_X2 FILLER_63_311 ();
 FILLCELL_X1 FILLER_63_313 ();
 FILLCELL_X4 FILLER_63_328 ();
 FILLCELL_X1 FILLER_63_332 ();
 FILLCELL_X8 FILLER_63_343 ();
 FILLCELL_X4 FILLER_63_351 ();
 FILLCELL_X2 FILLER_63_364 ();
 FILLCELL_X1 FILLER_63_366 ();
 FILLCELL_X4 FILLER_63_377 ();
 FILLCELL_X2 FILLER_63_381 ();
 FILLCELL_X4 FILLER_63_386 ();
 FILLCELL_X2 FILLER_63_390 ();
 FILLCELL_X2 FILLER_63_403 ();
 FILLCELL_X2 FILLER_63_416 ();
 FILLCELL_X16 FILLER_63_422 ();
 FILLCELL_X1 FILLER_63_438 ();
 FILLCELL_X1 FILLER_63_493 ();
 FILLCELL_X2 FILLER_63_507 ();
 FILLCELL_X2 FILLER_63_526 ();
 FILLCELL_X16 FILLER_63_533 ();
 FILLCELL_X2 FILLER_63_549 ();
 FILLCELL_X1 FILLER_63_551 ();
 FILLCELL_X2 FILLER_63_571 ();
 FILLCELL_X32 FILLER_63_607 ();
 FILLCELL_X16 FILLER_63_639 ();
 FILLCELL_X2 FILLER_63_663 ();
 FILLCELL_X1 FILLER_63_665 ();
 FILLCELL_X2 FILLER_63_670 ();
 FILLCELL_X1 FILLER_63_672 ();
 FILLCELL_X2 FILLER_63_681 ();
 FILLCELL_X8 FILLER_63_688 ();
 FILLCELL_X4 FILLER_63_706 ();
 FILLCELL_X16 FILLER_63_715 ();
 FILLCELL_X8 FILLER_63_731 ();
 FILLCELL_X2 FILLER_63_739 ();
 FILLCELL_X4 FILLER_63_756 ();
 FILLCELL_X8 FILLER_63_780 ();
 FILLCELL_X2 FILLER_63_788 ();
 FILLCELL_X1 FILLER_63_790 ();
 FILLCELL_X2 FILLER_63_802 ();
 FILLCELL_X1 FILLER_63_804 ();
 FILLCELL_X32 FILLER_63_822 ();
 FILLCELL_X8 FILLER_63_854 ();
 FILLCELL_X4 FILLER_63_862 ();
 FILLCELL_X2 FILLER_63_897 ();
 FILLCELL_X16 FILLER_63_911 ();
 FILLCELL_X4 FILLER_63_927 ();
 FILLCELL_X8 FILLER_63_941 ();
 FILLCELL_X2 FILLER_63_949 ();
 FILLCELL_X2 FILLER_63_957 ();
 FILLCELL_X2 FILLER_63_965 ();
 FILLCELL_X1 FILLER_63_967 ();
 FILLCELL_X2 FILLER_63_977 ();
 FILLCELL_X2 FILLER_63_986 ();
 FILLCELL_X4 FILLER_63_994 ();
 FILLCELL_X2 FILLER_63_998 ();
 FILLCELL_X16 FILLER_63_1009 ();
 FILLCELL_X2 FILLER_63_1025 ();
 FILLCELL_X2 FILLER_63_1040 ();
 FILLCELL_X1 FILLER_63_1098 ();
 FILLCELL_X2 FILLER_63_1114 ();
 FILLCELL_X1 FILLER_63_1116 ();
 FILLCELL_X16 FILLER_63_1121 ();
 FILLCELL_X1 FILLER_63_1137 ();
 FILLCELL_X4 FILLER_63_1163 ();
 FILLCELL_X1 FILLER_63_1167 ();
 FILLCELL_X2 FILLER_63_1175 ();
 FILLCELL_X8 FILLER_63_1194 ();
 FILLCELL_X4 FILLER_63_1202 ();
 FILLCELL_X2 FILLER_63_1206 ();
 FILLCELL_X1 FILLER_63_1208 ();
 FILLCELL_X32 FILLER_64_1 ();
 FILLCELL_X32 FILLER_64_33 ();
 FILLCELL_X8 FILLER_64_65 ();
 FILLCELL_X4 FILLER_64_73 ();
 FILLCELL_X2 FILLER_64_77 ();
 FILLCELL_X1 FILLER_64_79 ();
 FILLCELL_X16 FILLER_64_93 ();
 FILLCELL_X8 FILLER_64_109 ();
 FILLCELL_X2 FILLER_64_117 ();
 FILLCELL_X32 FILLER_64_132 ();
 FILLCELL_X32 FILLER_64_164 ();
 FILLCELL_X4 FILLER_64_196 ();
 FILLCELL_X2 FILLER_64_200 ();
 FILLCELL_X8 FILLER_64_215 ();
 FILLCELL_X4 FILLER_64_223 ();
 FILLCELL_X1 FILLER_64_227 ();
 FILLCELL_X4 FILLER_64_268 ();
 FILLCELL_X1 FILLER_64_272 ();
 FILLCELL_X2 FILLER_64_286 ();
 FILLCELL_X2 FILLER_64_301 ();
 FILLCELL_X1 FILLER_64_303 ();
 FILLCELL_X4 FILLER_64_339 ();
 FILLCELL_X1 FILLER_64_350 ();
 FILLCELL_X2 FILLER_64_358 ();
 FILLCELL_X1 FILLER_64_367 ();
 FILLCELL_X1 FILLER_64_373 ();
 FILLCELL_X8 FILLER_64_394 ();
 FILLCELL_X4 FILLER_64_402 ();
 FILLCELL_X1 FILLER_64_406 ();
 FILLCELL_X8 FILLER_64_425 ();
 FILLCELL_X4 FILLER_64_433 ();
 FILLCELL_X1 FILLER_64_437 ();
 FILLCELL_X16 FILLER_64_441 ();
 FILLCELL_X1 FILLER_64_457 ();
 FILLCELL_X2 FILLER_64_525 ();
 FILLCELL_X2 FILLER_64_534 ();
 FILLCELL_X2 FILLER_64_558 ();
 FILLCELL_X8 FILLER_64_581 ();
 FILLCELL_X16 FILLER_64_608 ();
 FILLCELL_X4 FILLER_64_624 ();
 FILLCELL_X2 FILLER_64_628 ();
 FILLCELL_X1 FILLER_64_630 ();
 FILLCELL_X8 FILLER_64_632 ();
 FILLCELL_X4 FILLER_64_640 ();
 FILLCELL_X2 FILLER_64_644 ();
 FILLCELL_X4 FILLER_64_649 ();
 FILLCELL_X2 FILLER_64_690 ();
 FILLCELL_X1 FILLER_64_692 ();
 FILLCELL_X2 FILLER_64_707 ();
 FILLCELL_X16 FILLER_64_712 ();
 FILLCELL_X2 FILLER_64_728 ();
 FILLCELL_X1 FILLER_64_730 ();
 FILLCELL_X1 FILLER_64_740 ();
 FILLCELL_X16 FILLER_64_745 ();
 FILLCELL_X1 FILLER_64_761 ();
 FILLCELL_X4 FILLER_64_765 ();
 FILLCELL_X8 FILLER_64_775 ();
 FILLCELL_X1 FILLER_64_783 ();
 FILLCELL_X4 FILLER_64_787 ();
 FILLCELL_X1 FILLER_64_791 ();
 FILLCELL_X2 FILLER_64_808 ();
 FILLCELL_X1 FILLER_64_810 ();
 FILLCELL_X32 FILLER_64_822 ();
 FILLCELL_X4 FILLER_64_854 ();
 FILLCELL_X2 FILLER_64_873 ();
 FILLCELL_X1 FILLER_64_875 ();
 FILLCELL_X2 FILLER_64_885 ();
 FILLCELL_X2 FILLER_64_928 ();
 FILLCELL_X1 FILLER_64_930 ();
 FILLCELL_X1 FILLER_64_947 ();
 FILLCELL_X8 FILLER_64_964 ();
 FILLCELL_X4 FILLER_64_972 ();
 FILLCELL_X4 FILLER_64_993 ();
 FILLCELL_X32 FILLER_64_1007 ();
 FILLCELL_X1 FILLER_64_1039 ();
 FILLCELL_X8 FILLER_64_1047 ();
 FILLCELL_X2 FILLER_64_1083 ();
 FILLCELL_X1 FILLER_64_1101 ();
 FILLCELL_X1 FILLER_64_1117 ();
 FILLCELL_X4 FILLER_64_1125 ();
 FILLCELL_X2 FILLER_64_1129 ();
 FILLCELL_X4 FILLER_64_1142 ();
 FILLCELL_X16 FILLER_64_1159 ();
 FILLCELL_X1 FILLER_64_1175 ();
 FILLCELL_X2 FILLER_64_1196 ();
 FILLCELL_X1 FILLER_64_1198 ();
 FILLCELL_X1 FILLER_64_1202 ();
 FILLCELL_X2 FILLER_64_1206 ();
 FILLCELL_X1 FILLER_64_1208 ();
 FILLCELL_X32 FILLER_65_1 ();
 FILLCELL_X32 FILLER_65_33 ();
 FILLCELL_X8 FILLER_65_65 ();
 FILLCELL_X4 FILLER_65_73 ();
 FILLCELL_X1 FILLER_65_77 ();
 FILLCELL_X4 FILLER_65_85 ();
 FILLCELL_X2 FILLER_65_89 ();
 FILLCELL_X32 FILLER_65_101 ();
 FILLCELL_X32 FILLER_65_133 ();
 FILLCELL_X1 FILLER_65_165 ();
 FILLCELL_X16 FILLER_65_173 ();
 FILLCELL_X4 FILLER_65_189 ();
 FILLCELL_X2 FILLER_65_193 ();
 FILLCELL_X1 FILLER_65_195 ();
 FILLCELL_X32 FILLER_65_200 ();
 FILLCELL_X8 FILLER_65_232 ();
 FILLCELL_X2 FILLER_65_240 ();
 FILLCELL_X1 FILLER_65_242 ();
 FILLCELL_X4 FILLER_65_260 ();
 FILLCELL_X2 FILLER_65_264 ();
 FILLCELL_X2 FILLER_65_279 ();
 FILLCELL_X1 FILLER_65_281 ();
 FILLCELL_X2 FILLER_65_285 ();
 FILLCELL_X4 FILLER_65_292 ();
 FILLCELL_X1 FILLER_65_296 ();
 FILLCELL_X2 FILLER_65_306 ();
 FILLCELL_X16 FILLER_65_315 ();
 FILLCELL_X4 FILLER_65_331 ();
 FILLCELL_X1 FILLER_65_335 ();
 FILLCELL_X8 FILLER_65_345 ();
 FILLCELL_X1 FILLER_65_353 ();
 FILLCELL_X4 FILLER_65_364 ();
 FILLCELL_X8 FILLER_65_385 ();
 FILLCELL_X32 FILLER_65_398 ();
 FILLCELL_X16 FILLER_65_430 ();
 FILLCELL_X8 FILLER_65_446 ();
 FILLCELL_X2 FILLER_65_454 ();
 FILLCELL_X1 FILLER_65_456 ();
 FILLCELL_X2 FILLER_65_474 ();
 FILLCELL_X2 FILLER_65_483 ();
 FILLCELL_X4 FILLER_65_512 ();
 FILLCELL_X4 FILLER_65_540 ();
 FILLCELL_X2 FILLER_65_544 ();
 FILLCELL_X4 FILLER_65_558 ();
 FILLCELL_X2 FILLER_65_562 ();
 FILLCELL_X1 FILLER_65_564 ();
 FILLCELL_X32 FILLER_65_576 ();
 FILLCELL_X16 FILLER_65_608 ();
 FILLCELL_X2 FILLER_65_624 ();
 FILLCELL_X1 FILLER_65_626 ();
 FILLCELL_X2 FILLER_65_654 ();
 FILLCELL_X1 FILLER_65_656 ();
 FILLCELL_X2 FILLER_65_678 ();
 FILLCELL_X1 FILLER_65_680 ();
 FILLCELL_X4 FILLER_65_701 ();
 FILLCELL_X4 FILLER_65_717 ();
 FILLCELL_X1 FILLER_65_721 ();
 FILLCELL_X1 FILLER_65_725 ();
 FILLCELL_X4 FILLER_65_744 ();
 FILLCELL_X2 FILLER_65_763 ();
 FILLCELL_X2 FILLER_65_772 ();
 FILLCELL_X1 FILLER_65_774 ();
 FILLCELL_X2 FILLER_65_782 ();
 FILLCELL_X16 FILLER_65_824 ();
 FILLCELL_X8 FILLER_65_840 ();
 FILLCELL_X4 FILLER_65_848 ();
 FILLCELL_X2 FILLER_65_852 ();
 FILLCELL_X1 FILLER_65_854 ();
 FILLCELL_X2 FILLER_65_876 ();
 FILLCELL_X1 FILLER_65_878 ();
 FILLCELL_X4 FILLER_65_889 ();
 FILLCELL_X1 FILLER_65_893 ();
 FILLCELL_X2 FILLER_65_932 ();
 FILLCELL_X2 FILLER_65_940 ();
 FILLCELL_X1 FILLER_65_942 ();
 FILLCELL_X4 FILLER_65_953 ();
 FILLCELL_X2 FILLER_65_957 ();
 FILLCELL_X1 FILLER_65_959 ();
 FILLCELL_X8 FILLER_65_978 ();
 FILLCELL_X1 FILLER_65_986 ();
 FILLCELL_X1 FILLER_65_996 ();
 FILLCELL_X2 FILLER_65_1015 ();
 FILLCELL_X1 FILLER_65_1017 ();
 FILLCELL_X2 FILLER_65_1027 ();
 FILLCELL_X2 FILLER_65_1043 ();
 FILLCELL_X1 FILLER_65_1045 ();
 FILLCELL_X4 FILLER_65_1060 ();
 FILLCELL_X2 FILLER_65_1064 ();
 FILLCELL_X1 FILLER_65_1099 ();
 FILLCELL_X2 FILLER_65_1109 ();
 FILLCELL_X1 FILLER_65_1111 ();
 FILLCELL_X8 FILLER_65_1129 ();
 FILLCELL_X4 FILLER_65_1137 ();
 FILLCELL_X2 FILLER_65_1141 ();
 FILLCELL_X2 FILLER_65_1149 ();
 FILLCELL_X1 FILLER_65_1151 ();
 FILLCELL_X1 FILLER_65_1156 ();
 FILLCELL_X4 FILLER_65_1172 ();
 FILLCELL_X2 FILLER_65_1176 ();
 FILLCELL_X1 FILLER_65_1178 ();
 FILLCELL_X8 FILLER_65_1201 ();
 FILLCELL_X16 FILLER_66_1 ();
 FILLCELL_X8 FILLER_66_17 ();
 FILLCELL_X2 FILLER_66_25 ();
 FILLCELL_X4 FILLER_66_30 ();
 FILLCELL_X2 FILLER_66_34 ();
 FILLCELL_X16 FILLER_66_65 ();
 FILLCELL_X2 FILLER_66_98 ();
 FILLCELL_X1 FILLER_66_100 ();
 FILLCELL_X8 FILLER_66_108 ();
 FILLCELL_X2 FILLER_66_116 ();
 FILLCELL_X1 FILLER_66_118 ();
 FILLCELL_X1 FILLER_66_132 ();
 FILLCELL_X8 FILLER_66_147 ();
 FILLCELL_X2 FILLER_66_155 ();
 FILLCELL_X2 FILLER_66_181 ();
 FILLCELL_X4 FILLER_66_197 ();
 FILLCELL_X2 FILLER_66_208 ();
 FILLCELL_X1 FILLER_66_217 ();
 FILLCELL_X32 FILLER_66_253 ();
 FILLCELL_X2 FILLER_66_285 ();
 FILLCELL_X1 FILLER_66_287 ();
 FILLCELL_X2 FILLER_66_292 ();
 FILLCELL_X1 FILLER_66_294 ();
 FILLCELL_X4 FILLER_66_312 ();
 FILLCELL_X1 FILLER_66_342 ();
 FILLCELL_X4 FILLER_66_377 ();
 FILLCELL_X1 FILLER_66_381 ();
 FILLCELL_X16 FILLER_66_400 ();
 FILLCELL_X2 FILLER_66_416 ();
 FILLCELL_X1 FILLER_66_431 ();
 FILLCELL_X4 FILLER_66_448 ();
 FILLCELL_X1 FILLER_66_455 ();
 FILLCELL_X1 FILLER_66_478 ();
 FILLCELL_X2 FILLER_66_510 ();
 FILLCELL_X1 FILLER_66_551 ();
 FILLCELL_X1 FILLER_66_562 ();
 FILLCELL_X1 FILLER_66_587 ();
 FILLCELL_X8 FILLER_66_596 ();
 FILLCELL_X2 FILLER_66_604 ();
 FILLCELL_X8 FILLER_66_632 ();
 FILLCELL_X4 FILLER_66_640 ();
 FILLCELL_X1 FILLER_66_644 ();
 FILLCELL_X1 FILLER_66_664 ();
 FILLCELL_X8 FILLER_66_668 ();
 FILLCELL_X1 FILLER_66_676 ();
 FILLCELL_X8 FILLER_66_690 ();
 FILLCELL_X4 FILLER_66_698 ();
 FILLCELL_X1 FILLER_66_702 ();
 FILLCELL_X2 FILLER_66_710 ();
 FILLCELL_X8 FILLER_66_719 ();
 FILLCELL_X4 FILLER_66_727 ();
 FILLCELL_X2 FILLER_66_731 ();
 FILLCELL_X1 FILLER_66_733 ();
 FILLCELL_X8 FILLER_66_743 ();
 FILLCELL_X2 FILLER_66_751 ();
 FILLCELL_X1 FILLER_66_753 ();
 FILLCELL_X1 FILLER_66_768 ();
 FILLCELL_X8 FILLER_66_773 ();
 FILLCELL_X2 FILLER_66_781 ();
 FILLCELL_X1 FILLER_66_783 ();
 FILLCELL_X1 FILLER_66_797 ();
 FILLCELL_X32 FILLER_66_821 ();
 FILLCELL_X4 FILLER_66_853 ();
 FILLCELL_X1 FILLER_66_877 ();
 FILLCELL_X1 FILLER_66_891 ();
 FILLCELL_X2 FILLER_66_906 ();
 FILLCELL_X2 FILLER_66_912 ();
 FILLCELL_X4 FILLER_66_920 ();
 FILLCELL_X2 FILLER_66_924 ();
 FILLCELL_X1 FILLER_66_926 ();
 FILLCELL_X1 FILLER_66_940 ();
 FILLCELL_X4 FILLER_66_951 ();
 FILLCELL_X2 FILLER_66_965 ();
 FILLCELL_X1 FILLER_66_967 ();
 FILLCELL_X4 FILLER_66_1001 ();
 FILLCELL_X1 FILLER_66_1005 ();
 FILLCELL_X8 FILLER_66_1013 ();
 FILLCELL_X2 FILLER_66_1021 ();
 FILLCELL_X4 FILLER_66_1046 ();
 FILLCELL_X1 FILLER_66_1050 ();
 FILLCELL_X2 FILLER_66_1064 ();
 FILLCELL_X1 FILLER_66_1066 ();
 FILLCELL_X4 FILLER_66_1078 ();
 FILLCELL_X2 FILLER_66_1096 ();
 FILLCELL_X1 FILLER_66_1098 ();
 FILLCELL_X4 FILLER_66_1103 ();
 FILLCELL_X2 FILLER_66_1107 ();
 FILLCELL_X1 FILLER_66_1109 ();
 FILLCELL_X1 FILLER_66_1117 ();
 FILLCELL_X8 FILLER_66_1124 ();
 FILLCELL_X2 FILLER_66_1132 ();
 FILLCELL_X1 FILLER_66_1134 ();
 FILLCELL_X2 FILLER_66_1146 ();
 FILLCELL_X4 FILLER_66_1160 ();
 FILLCELL_X2 FILLER_66_1164 ();
 FILLCELL_X1 FILLER_66_1166 ();
 FILLCELL_X4 FILLER_66_1180 ();
 FILLCELL_X4 FILLER_66_1199 ();
 FILLCELL_X16 FILLER_67_1 ();
 FILLCELL_X8 FILLER_67_17 ();
 FILLCELL_X2 FILLER_67_25 ();
 FILLCELL_X16 FILLER_67_53 ();
 FILLCELL_X4 FILLER_67_69 ();
 FILLCELL_X8 FILLER_67_94 ();
 FILLCELL_X4 FILLER_67_102 ();
 FILLCELL_X2 FILLER_67_126 ();
 FILLCELL_X2 FILLER_67_131 ();
 FILLCELL_X16 FILLER_67_158 ();
 FILLCELL_X4 FILLER_67_174 ();
 FILLCELL_X2 FILLER_67_178 ();
 FILLCELL_X1 FILLER_67_180 ();
 FILLCELL_X2 FILLER_67_209 ();
 FILLCELL_X1 FILLER_67_211 ();
 FILLCELL_X2 FILLER_67_239 ();
 FILLCELL_X16 FILLER_67_244 ();
 FILLCELL_X4 FILLER_67_260 ();
 FILLCELL_X2 FILLER_67_264 ();
 FILLCELL_X4 FILLER_67_273 ();
 FILLCELL_X4 FILLER_67_280 ();
 FILLCELL_X2 FILLER_67_310 ();
 FILLCELL_X1 FILLER_67_312 ();
 FILLCELL_X16 FILLER_67_318 ();
 FILLCELL_X8 FILLER_67_334 ();
 FILLCELL_X2 FILLER_67_342 ();
 FILLCELL_X4 FILLER_67_347 ();
 FILLCELL_X2 FILLER_67_351 ();
 FILLCELL_X8 FILLER_67_355 ();
 FILLCELL_X4 FILLER_67_363 ();
 FILLCELL_X2 FILLER_67_367 ();
 FILLCELL_X1 FILLER_67_471 ();
 FILLCELL_X1 FILLER_67_491 ();
 FILLCELL_X1 FILLER_67_496 ();
 FILLCELL_X8 FILLER_67_527 ();
 FILLCELL_X2 FILLER_67_535 ();
 FILLCELL_X8 FILLER_67_572 ();
 FILLCELL_X4 FILLER_67_580 ();
 FILLCELL_X2 FILLER_67_590 ();
 FILLCELL_X1 FILLER_67_596 ();
 FILLCELL_X32 FILLER_67_601 ();
 FILLCELL_X8 FILLER_67_633 ();
 FILLCELL_X2 FILLER_67_641 ();
 FILLCELL_X1 FILLER_67_655 ();
 FILLCELL_X8 FILLER_67_671 ();
 FILLCELL_X2 FILLER_67_679 ();
 FILLCELL_X2 FILLER_67_694 ();
 FILLCELL_X1 FILLER_67_703 ();
 FILLCELL_X8 FILLER_67_718 ();
 FILLCELL_X4 FILLER_67_726 ();
 FILLCELL_X1 FILLER_67_730 ();
 FILLCELL_X1 FILLER_67_743 ();
 FILLCELL_X2 FILLER_67_751 ();
 FILLCELL_X1 FILLER_67_764 ();
 FILLCELL_X1 FILLER_67_771 ();
 FILLCELL_X16 FILLER_67_778 ();
 FILLCELL_X8 FILLER_67_794 ();
 FILLCELL_X2 FILLER_67_802 ();
 FILLCELL_X1 FILLER_67_804 ();
 FILLCELL_X32 FILLER_67_828 ();
 FILLCELL_X2 FILLER_67_860 ();
 FILLCELL_X1 FILLER_67_866 ();
 FILLCELL_X2 FILLER_67_879 ();
 FILLCELL_X2 FILLER_67_890 ();
 FILLCELL_X1 FILLER_67_892 ();
 FILLCELL_X1 FILLER_67_902 ();
 FILLCELL_X2 FILLER_67_910 ();
 FILLCELL_X2 FILLER_67_924 ();
 FILLCELL_X1 FILLER_67_926 ();
 FILLCELL_X1 FILLER_67_952 ();
 FILLCELL_X16 FILLER_67_977 ();
 FILLCELL_X1 FILLER_67_993 ();
 FILLCELL_X16 FILLER_67_1011 ();
 FILLCELL_X1 FILLER_67_1032 ();
 FILLCELL_X2 FILLER_67_1047 ();
 FILLCELL_X1 FILLER_67_1049 ();
 FILLCELL_X1 FILLER_67_1063 ();
 FILLCELL_X2 FILLER_67_1069 ();
 FILLCELL_X1 FILLER_67_1071 ();
 FILLCELL_X2 FILLER_67_1085 ();
 FILLCELL_X1 FILLER_67_1098 ();
 FILLCELL_X4 FILLER_67_1110 ();
 FILLCELL_X1 FILLER_67_1114 ();
 FILLCELL_X8 FILLER_67_1124 ();
 FILLCELL_X2 FILLER_67_1132 ();
 FILLCELL_X1 FILLER_67_1134 ();
 FILLCELL_X4 FILLER_67_1141 ();
 FILLCELL_X2 FILLER_67_1145 ();
 FILLCELL_X1 FILLER_67_1147 ();
 FILLCELL_X2 FILLER_67_1160 ();
 FILLCELL_X1 FILLER_67_1162 ();
 FILLCELL_X4 FILLER_67_1171 ();
 FILLCELL_X2 FILLER_67_1175 ();
 FILLCELL_X1 FILLER_67_1177 ();
 FILLCELL_X2 FILLER_67_1203 ();
 FILLCELL_X16 FILLER_68_4 ();
 FILLCELL_X2 FILLER_68_20 ();
 FILLCELL_X1 FILLER_68_22 ();
 FILLCELL_X16 FILLER_68_49 ();
 FILLCELL_X8 FILLER_68_65 ();
 FILLCELL_X1 FILLER_68_117 ();
 FILLCELL_X2 FILLER_68_189 ();
 FILLCELL_X1 FILLER_68_198 ();
 FILLCELL_X4 FILLER_68_206 ();
 FILLCELL_X1 FILLER_68_224 ();
 FILLCELL_X2 FILLER_68_250 ();
 FILLCELL_X1 FILLER_68_252 ();
 FILLCELL_X1 FILLER_68_273 ();
 FILLCELL_X4 FILLER_68_290 ();
 FILLCELL_X2 FILLER_68_294 ();
 FILLCELL_X1 FILLER_68_310 ();
 FILLCELL_X4 FILLER_68_324 ();
 FILLCELL_X8 FILLER_68_331 ();
 FILLCELL_X4 FILLER_68_339 ();
 FILLCELL_X2 FILLER_68_358 ();
 FILLCELL_X1 FILLER_68_360 ();
 FILLCELL_X2 FILLER_68_364 ();
 FILLCELL_X1 FILLER_68_366 ();
 FILLCELL_X2 FILLER_68_390 ();
 FILLCELL_X8 FILLER_68_407 ();
 FILLCELL_X1 FILLER_68_497 ();
 FILLCELL_X4 FILLER_68_513 ();
 FILLCELL_X1 FILLER_68_517 ();
 FILLCELL_X8 FILLER_68_579 ();
 FILLCELL_X2 FILLER_68_591 ();
 FILLCELL_X1 FILLER_68_593 ();
 FILLCELL_X2 FILLER_68_597 ();
 FILLCELL_X16 FILLER_68_610 ();
 FILLCELL_X4 FILLER_68_626 ();
 FILLCELL_X1 FILLER_68_630 ();
 FILLCELL_X4 FILLER_68_632 ();
 FILLCELL_X1 FILLER_68_636 ();
 FILLCELL_X4 FILLER_68_648 ();
 FILLCELL_X4 FILLER_68_655 ();
 FILLCELL_X16 FILLER_68_665 ();
 FILLCELL_X4 FILLER_68_681 ();
 FILLCELL_X1 FILLER_68_685 ();
 FILLCELL_X4 FILLER_68_690 ();
 FILLCELL_X1 FILLER_68_694 ();
 FILLCELL_X8 FILLER_68_710 ();
 FILLCELL_X4 FILLER_68_718 ();
 FILLCELL_X2 FILLER_68_722 ();
 FILLCELL_X4 FILLER_68_727 ();
 FILLCELL_X2 FILLER_68_731 ();
 FILLCELL_X4 FILLER_68_737 ();
 FILLCELL_X2 FILLER_68_741 ();
 FILLCELL_X16 FILLER_68_747 ();
 FILLCELL_X1 FILLER_68_763 ();
 FILLCELL_X2 FILLER_68_771 ();
 FILLCELL_X2 FILLER_68_793 ();
 FILLCELL_X1 FILLER_68_800 ();
 FILLCELL_X2 FILLER_68_805 ();
 FILLCELL_X1 FILLER_68_807 ();
 FILLCELL_X8 FILLER_68_820 ();
 FILLCELL_X2 FILLER_68_828 ();
 FILLCELL_X16 FILLER_68_840 ();
 FILLCELL_X8 FILLER_68_856 ();
 FILLCELL_X8 FILLER_68_873 ();
 FILLCELL_X4 FILLER_68_881 ();
 FILLCELL_X1 FILLER_68_895 ();
 FILLCELL_X2 FILLER_68_929 ();
 FILLCELL_X8 FILLER_68_944 ();
 FILLCELL_X2 FILLER_68_952 ();
 FILLCELL_X1 FILLER_68_954 ();
 FILLCELL_X2 FILLER_68_969 ();
 FILLCELL_X1 FILLER_68_981 ();
 FILLCELL_X16 FILLER_68_989 ();
 FILLCELL_X1 FILLER_68_1005 ();
 FILLCELL_X2 FILLER_68_1023 ();
 FILLCELL_X1 FILLER_68_1025 ();
 FILLCELL_X4 FILLER_68_1035 ();
 FILLCELL_X1 FILLER_68_1059 ();
 FILLCELL_X4 FILLER_68_1074 ();
 FILLCELL_X1 FILLER_68_1078 ();
 FILLCELL_X4 FILLER_68_1083 ();
 FILLCELL_X4 FILLER_68_1096 ();
 FILLCELL_X2 FILLER_68_1100 ();
 FILLCELL_X1 FILLER_68_1119 ();
 FILLCELL_X1 FILLER_68_1123 ();
 FILLCELL_X2 FILLER_68_1154 ();
 FILLCELL_X8 FILLER_68_1169 ();
 FILLCELL_X4 FILLER_68_1177 ();
 FILLCELL_X2 FILLER_68_1181 ();
 FILLCELL_X1 FILLER_68_1200 ();
 FILLCELL_X4 FILLER_68_1204 ();
 FILLCELL_X1 FILLER_68_1208 ();
 FILLCELL_X16 FILLER_69_1 ();
 FILLCELL_X4 FILLER_69_17 ();
 FILLCELL_X2 FILLER_69_21 ();
 FILLCELL_X8 FILLER_69_27 ();
 FILLCELL_X4 FILLER_69_35 ();
 FILLCELL_X2 FILLER_69_39 ();
 FILLCELL_X1 FILLER_69_41 ();
 FILLCELL_X16 FILLER_69_49 ();
 FILLCELL_X8 FILLER_69_65 ();
 FILLCELL_X4 FILLER_69_73 ();
 FILLCELL_X8 FILLER_69_87 ();
 FILLCELL_X4 FILLER_69_95 ();
 FILLCELL_X2 FILLER_69_99 ();
 FILLCELL_X4 FILLER_69_111 ();
 FILLCELL_X1 FILLER_69_148 ();
 FILLCELL_X4 FILLER_69_157 ();
 FILLCELL_X1 FILLER_69_182 ();
 FILLCELL_X1 FILLER_69_194 ();
 FILLCELL_X2 FILLER_69_201 ();
 FILLCELL_X1 FILLER_69_203 ();
 FILLCELL_X2 FILLER_69_229 ();
 FILLCELL_X2 FILLER_69_251 ();
 FILLCELL_X1 FILLER_69_253 ();
 FILLCELL_X16 FILLER_69_263 ();
 FILLCELL_X4 FILLER_69_279 ();
 FILLCELL_X4 FILLER_69_290 ();
 FILLCELL_X1 FILLER_69_311 ();
 FILLCELL_X2 FILLER_69_319 ();
 FILLCELL_X2 FILLER_69_325 ();
 FILLCELL_X8 FILLER_69_336 ();
 FILLCELL_X2 FILLER_69_344 ();
 FILLCELL_X1 FILLER_69_346 ();
 FILLCELL_X16 FILLER_69_356 ();
 FILLCELL_X2 FILLER_69_394 ();
 FILLCELL_X1 FILLER_69_396 ();
 FILLCELL_X8 FILLER_69_410 ();
 FILLCELL_X4 FILLER_69_418 ();
 FILLCELL_X2 FILLER_69_422 ();
 FILLCELL_X1 FILLER_69_424 ();
 FILLCELL_X8 FILLER_69_438 ();
 FILLCELL_X4 FILLER_69_507 ();
 FILLCELL_X1 FILLER_69_511 ();
 FILLCELL_X2 FILLER_69_515 ();
 FILLCELL_X1 FILLER_69_517 ();
 FILLCELL_X2 FILLER_69_527 ();
 FILLCELL_X1 FILLER_69_529 ();
 FILLCELL_X2 FILLER_69_536 ();
 FILLCELL_X8 FILLER_69_569 ();
 FILLCELL_X4 FILLER_69_577 ();
 FILLCELL_X2 FILLER_69_581 ();
 FILLCELL_X1 FILLER_69_583 ();
 FILLCELL_X32 FILLER_69_601 ();
 FILLCELL_X8 FILLER_69_633 ();
 FILLCELL_X4 FILLER_69_641 ();
 FILLCELL_X2 FILLER_69_660 ();
 FILLCELL_X1 FILLER_69_662 ();
 FILLCELL_X8 FILLER_69_666 ();
 FILLCELL_X2 FILLER_69_674 ();
 FILLCELL_X1 FILLER_69_676 ();
 FILLCELL_X1 FILLER_69_691 ();
 FILLCELL_X2 FILLER_69_701 ();
 FILLCELL_X1 FILLER_69_703 ();
 FILLCELL_X4 FILLER_69_718 ();
 FILLCELL_X2 FILLER_69_722 ();
 FILLCELL_X2 FILLER_69_731 ();
 FILLCELL_X1 FILLER_69_758 ();
 FILLCELL_X16 FILLER_69_766 ();
 FILLCELL_X4 FILLER_69_782 ();
 FILLCELL_X2 FILLER_69_802 ();
 FILLCELL_X8 FILLER_69_827 ();
 FILLCELL_X8 FILLER_69_844 ();
 FILLCELL_X2 FILLER_69_852 ();
 FILLCELL_X1 FILLER_69_854 ();
 FILLCELL_X4 FILLER_69_858 ();
 FILLCELL_X2 FILLER_69_862 ();
 FILLCELL_X1 FILLER_69_864 ();
 FILLCELL_X16 FILLER_69_879 ();
 FILLCELL_X4 FILLER_69_895 ();
 FILLCELL_X2 FILLER_69_908 ();
 FILLCELL_X2 FILLER_69_916 ();
 FILLCELL_X4 FILLER_69_941 ();
 FILLCELL_X2 FILLER_69_945 ();
 FILLCELL_X1 FILLER_69_947 ();
 FILLCELL_X8 FILLER_69_974 ();
 FILLCELL_X8 FILLER_69_989 ();
 FILLCELL_X2 FILLER_69_1012 ();
 FILLCELL_X1 FILLER_69_1014 ();
 FILLCELL_X16 FILLER_69_1019 ();
 FILLCELL_X1 FILLER_69_1035 ();
 FILLCELL_X4 FILLER_69_1045 ();
 FILLCELL_X4 FILLER_69_1063 ();
 FILLCELL_X8 FILLER_69_1071 ();
 FILLCELL_X4 FILLER_69_1079 ();
 FILLCELL_X1 FILLER_69_1083 ();
 FILLCELL_X4 FILLER_69_1087 ();
 FILLCELL_X8 FILLER_69_1102 ();
 FILLCELL_X2 FILLER_69_1110 ();
 FILLCELL_X1 FILLER_69_1112 ();
 FILLCELL_X2 FILLER_69_1117 ();
 FILLCELL_X4 FILLER_69_1126 ();
 FILLCELL_X2 FILLER_69_1130 ();
 FILLCELL_X1 FILLER_69_1132 ();
 FILLCELL_X8 FILLER_69_1138 ();
 FILLCELL_X4 FILLER_69_1146 ();
 FILLCELL_X16 FILLER_69_1180 ();
 FILLCELL_X4 FILLER_69_1196 ();
 FILLCELL_X1 FILLER_69_1200 ();
 FILLCELL_X1 FILLER_69_1204 ();
 FILLCELL_X32 FILLER_70_1 ();
 FILLCELL_X8 FILLER_70_33 ();
 FILLCELL_X2 FILLER_70_41 ();
 FILLCELL_X16 FILLER_70_62 ();
 FILLCELL_X8 FILLER_70_78 ();
 FILLCELL_X4 FILLER_70_105 ();
 FILLCELL_X2 FILLER_70_109 ();
 FILLCELL_X1 FILLER_70_111 ();
 FILLCELL_X8 FILLER_70_116 ();
 FILLCELL_X2 FILLER_70_128 ();
 FILLCELL_X1 FILLER_70_130 ();
 FILLCELL_X2 FILLER_70_135 ();
 FILLCELL_X1 FILLER_70_148 ();
 FILLCELL_X4 FILLER_70_153 ();
 FILLCELL_X2 FILLER_70_157 ();
 FILLCELL_X1 FILLER_70_159 ();
 FILLCELL_X4 FILLER_70_167 ();
 FILLCELL_X4 FILLER_70_198 ();
 FILLCELL_X2 FILLER_70_202 ();
 FILLCELL_X2 FILLER_70_222 ();
 FILLCELL_X1 FILLER_70_231 ();
 FILLCELL_X8 FILLER_70_252 ();
 FILLCELL_X4 FILLER_70_260 ();
 FILLCELL_X1 FILLER_70_264 ();
 FILLCELL_X4 FILLER_70_282 ();
 FILLCELL_X2 FILLER_70_286 ();
 FILLCELL_X1 FILLER_70_288 ();
 FILLCELL_X1 FILLER_70_292 ();
 FILLCELL_X2 FILLER_70_297 ();
 FILLCELL_X1 FILLER_70_299 ();
 FILLCELL_X1 FILLER_70_313 ();
 FILLCELL_X8 FILLER_70_318 ();
 FILLCELL_X2 FILLER_70_326 ();
 FILLCELL_X2 FILLER_70_331 ();
 FILLCELL_X16 FILLER_70_353 ();
 FILLCELL_X1 FILLER_70_369 ();
 FILLCELL_X16 FILLER_70_399 ();
 FILLCELL_X4 FILLER_70_415 ();
 FILLCELL_X2 FILLER_70_419 ();
 FILLCELL_X1 FILLER_70_421 ();
 FILLCELL_X4 FILLER_70_448 ();
 FILLCELL_X1 FILLER_70_452 ();
 FILLCELL_X2 FILLER_70_462 ();
 FILLCELL_X8 FILLER_70_509 ();
 FILLCELL_X1 FILLER_70_517 ();
 FILLCELL_X1 FILLER_70_528 ();
 FILLCELL_X4 FILLER_70_535 ();
 FILLCELL_X4 FILLER_70_543 ();
 FILLCELL_X2 FILLER_70_547 ();
 FILLCELL_X2 FILLER_70_587 ();
 FILLCELL_X1 FILLER_70_589 ();
 FILLCELL_X16 FILLER_70_614 ();
 FILLCELL_X1 FILLER_70_630 ();
 FILLCELL_X8 FILLER_70_632 ();
 FILLCELL_X4 FILLER_70_640 ();
 FILLCELL_X2 FILLER_70_644 ();
 FILLCELL_X16 FILLER_70_652 ();
 FILLCELL_X8 FILLER_70_688 ();
 FILLCELL_X1 FILLER_70_704 ();
 FILLCELL_X2 FILLER_70_724 ();
 FILLCELL_X1 FILLER_70_732 ();
 FILLCELL_X2 FILLER_70_738 ();
 FILLCELL_X4 FILLER_70_758 ();
 FILLCELL_X2 FILLER_70_762 ();
 FILLCELL_X1 FILLER_70_780 ();
 FILLCELL_X2 FILLER_70_785 ();
 FILLCELL_X2 FILLER_70_791 ();
 FILLCELL_X2 FILLER_70_807 ();
 FILLCELL_X8 FILLER_70_838 ();
 FILLCELL_X4 FILLER_70_846 ();
 FILLCELL_X2 FILLER_70_886 ();
 FILLCELL_X1 FILLER_70_895 ();
 FILLCELL_X2 FILLER_70_911 ();
 FILLCELL_X1 FILLER_70_913 ();
 FILLCELL_X4 FILLER_70_916 ();
 FILLCELL_X1 FILLER_70_920 ();
 FILLCELL_X16 FILLER_70_948 ();
 FILLCELL_X8 FILLER_70_964 ();
 FILLCELL_X2 FILLER_70_972 ();
 FILLCELL_X2 FILLER_70_980 ();
 FILLCELL_X4 FILLER_70_994 ();
 FILLCELL_X2 FILLER_70_998 ();
 FILLCELL_X1 FILLER_70_1000 ();
 FILLCELL_X4 FILLER_70_1011 ();
 FILLCELL_X2 FILLER_70_1015 ();
 FILLCELL_X1 FILLER_70_1017 ();
 FILLCELL_X2 FILLER_70_1031 ();
 FILLCELL_X16 FILLER_70_1036 ();
 FILLCELL_X4 FILLER_70_1063 ();
 FILLCELL_X2 FILLER_70_1067 ();
 FILLCELL_X1 FILLER_70_1069 ();
 FILLCELL_X8 FILLER_70_1084 ();
 FILLCELL_X1 FILLER_70_1092 ();
 FILLCELL_X1 FILLER_70_1105 ();
 FILLCELL_X1 FILLER_70_1110 ();
 FILLCELL_X4 FILLER_70_1116 ();
 FILLCELL_X2 FILLER_70_1120 ();
 FILLCELL_X2 FILLER_70_1133 ();
 FILLCELL_X1 FILLER_70_1135 ();
 FILLCELL_X16 FILLER_70_1140 ();
 FILLCELL_X4 FILLER_70_1156 ();
 FILLCELL_X2 FILLER_70_1167 ();
 FILLCELL_X4 FILLER_70_1180 ();
 FILLCELL_X1 FILLER_70_1184 ();
 FILLCELL_X16 FILLER_70_1192 ();
 FILLCELL_X1 FILLER_70_1208 ();
 FILLCELL_X4 FILLER_71_1 ();
 FILLCELL_X8 FILLER_71_9 ();
 FILLCELL_X2 FILLER_71_17 ();
 FILLCELL_X1 FILLER_71_19 ();
 FILLCELL_X4 FILLER_71_30 ();
 FILLCELL_X16 FILLER_71_51 ();
 FILLCELL_X8 FILLER_71_67 ();
 FILLCELL_X4 FILLER_71_75 ();
 FILLCELL_X2 FILLER_71_79 ();
 FILLCELL_X1 FILLER_71_95 ();
 FILLCELL_X2 FILLER_71_109 ();
 FILLCELL_X1 FILLER_71_114 ();
 FILLCELL_X1 FILLER_71_121 ();
 FILLCELL_X2 FILLER_71_126 ();
 FILLCELL_X2 FILLER_71_136 ();
 FILLCELL_X1 FILLER_71_138 ();
 FILLCELL_X8 FILLER_71_158 ();
 FILLCELL_X1 FILLER_71_183 ();
 FILLCELL_X8 FILLER_71_197 ();
 FILLCELL_X1 FILLER_71_205 ();
 FILLCELL_X1 FILLER_71_215 ();
 FILLCELL_X1 FILLER_71_227 ();
 FILLCELL_X1 FILLER_71_238 ();
 FILLCELL_X4 FILLER_71_246 ();
 FILLCELL_X1 FILLER_71_250 ();
 FILLCELL_X32 FILLER_71_258 ();
 FILLCELL_X2 FILLER_71_290 ();
 FILLCELL_X4 FILLER_71_301 ();
 FILLCELL_X2 FILLER_71_305 ();
 FILLCELL_X1 FILLER_71_307 ();
 FILLCELL_X8 FILLER_71_315 ();
 FILLCELL_X4 FILLER_71_323 ();
 FILLCELL_X2 FILLER_71_327 ();
 FILLCELL_X4 FILLER_71_349 ();
 FILLCELL_X2 FILLER_71_375 ();
 FILLCELL_X4 FILLER_71_389 ();
 FILLCELL_X1 FILLER_71_393 ();
 FILLCELL_X4 FILLER_71_401 ();
 FILLCELL_X1 FILLER_71_405 ();
 FILLCELL_X16 FILLER_71_420 ();
 FILLCELL_X8 FILLER_71_436 ();
 FILLCELL_X2 FILLER_71_444 ();
 FILLCELL_X1 FILLER_71_446 ();
 FILLCELL_X4 FILLER_71_460 ();
 FILLCELL_X1 FILLER_71_495 ();
 FILLCELL_X1 FILLER_71_534 ();
 FILLCELL_X2 FILLER_71_581 ();
 FILLCELL_X1 FILLER_71_583 ();
 FILLCELL_X32 FILLER_71_600 ();
 FILLCELL_X16 FILLER_71_632 ();
 FILLCELL_X2 FILLER_71_648 ();
 FILLCELL_X4 FILLER_71_657 ();
 FILLCELL_X1 FILLER_71_661 ();
 FILLCELL_X2 FILLER_71_665 ();
 FILLCELL_X8 FILLER_71_700 ();
 FILLCELL_X1 FILLER_71_708 ();
 FILLCELL_X1 FILLER_71_744 ();
 FILLCELL_X1 FILLER_71_782 ();
 FILLCELL_X2 FILLER_71_801 ();
 FILLCELL_X2 FILLER_71_816 ();
 FILLCELL_X32 FILLER_71_831 ();
 FILLCELL_X8 FILLER_71_869 ();
 FILLCELL_X4 FILLER_71_877 ();
 FILLCELL_X2 FILLER_71_881 ();
 FILLCELL_X2 FILLER_71_893 ();
 FILLCELL_X1 FILLER_71_934 ();
 FILLCELL_X2 FILLER_71_959 ();
 FILLCELL_X2 FILLER_71_968 ();
 FILLCELL_X1 FILLER_71_970 ();
 FILLCELL_X16 FILLER_71_992 ();
 FILLCELL_X4 FILLER_71_1008 ();
 FILLCELL_X1 FILLER_71_1012 ();
 FILLCELL_X4 FILLER_71_1022 ();
 FILLCELL_X2 FILLER_71_1026 ();
 FILLCELL_X1 FILLER_71_1028 ();
 FILLCELL_X4 FILLER_71_1072 ();
 FILLCELL_X2 FILLER_71_1076 ();
 FILLCELL_X4 FILLER_71_1082 ();
 FILLCELL_X4 FILLER_71_1100 ();
 FILLCELL_X1 FILLER_71_1104 ();
 FILLCELL_X4 FILLER_71_1118 ();
 FILLCELL_X2 FILLER_71_1122 ();
 FILLCELL_X8 FILLER_71_1128 ();
 FILLCELL_X4 FILLER_71_1142 ();
 FILLCELL_X2 FILLER_71_1146 ();
 FILLCELL_X1 FILLER_71_1148 ();
 FILLCELL_X2 FILLER_71_1156 ();
 FILLCELL_X1 FILLER_71_1158 ();
 FILLCELL_X1 FILLER_71_1166 ();
 FILLCELL_X16 FILLER_71_1178 ();
 FILLCELL_X8 FILLER_71_1197 ();
 FILLCELL_X4 FILLER_71_1205 ();
 FILLCELL_X16 FILLER_72_1 ();
 FILLCELL_X8 FILLER_72_17 ();
 FILLCELL_X8 FILLER_72_51 ();
 FILLCELL_X4 FILLER_72_59 ();
 FILLCELL_X2 FILLER_72_63 ();
 FILLCELL_X1 FILLER_72_65 ();
 FILLCELL_X1 FILLER_72_86 ();
 FILLCELL_X1 FILLER_72_94 ();
 FILLCELL_X1 FILLER_72_152 ();
 FILLCELL_X1 FILLER_72_157 ();
 FILLCELL_X2 FILLER_72_193 ();
 FILLCELL_X1 FILLER_72_195 ();
 FILLCELL_X2 FILLER_72_201 ();
 FILLCELL_X1 FILLER_72_203 ();
 FILLCELL_X2 FILLER_72_207 ();
 FILLCELL_X1 FILLER_72_209 ();
 FILLCELL_X1 FILLER_72_248 ();
 FILLCELL_X2 FILLER_72_254 ();
 FILLCELL_X1 FILLER_72_256 ();
 FILLCELL_X16 FILLER_72_264 ();
 FILLCELL_X1 FILLER_72_280 ();
 FILLCELL_X2 FILLER_72_286 ();
 FILLCELL_X1 FILLER_72_288 ();
 FILLCELL_X8 FILLER_72_306 ();
 FILLCELL_X4 FILLER_72_314 ();
 FILLCELL_X1 FILLER_72_318 ();
 FILLCELL_X1 FILLER_72_339 ();
 FILLCELL_X8 FILLER_72_357 ();
 FILLCELL_X2 FILLER_72_365 ();
 FILLCELL_X1 FILLER_72_367 ();
 FILLCELL_X16 FILLER_72_389 ();
 FILLCELL_X1 FILLER_72_405 ();
 FILLCELL_X8 FILLER_72_410 ();
 FILLCELL_X4 FILLER_72_418 ();
 FILLCELL_X1 FILLER_72_458 ();
 FILLCELL_X2 FILLER_72_469 ();
 FILLCELL_X2 FILLER_72_480 ();
 FILLCELL_X2 FILLER_72_485 ();
 FILLCELL_X8 FILLER_72_516 ();
 FILLCELL_X1 FILLER_72_524 ();
 FILLCELL_X4 FILLER_72_535 ();
 FILLCELL_X1 FILLER_72_539 ();
 FILLCELL_X2 FILLER_72_564 ();
 FILLCELL_X1 FILLER_72_566 ();
 FILLCELL_X4 FILLER_72_581 ();
 FILLCELL_X1 FILLER_72_585 ();
 FILLCELL_X4 FILLER_72_615 ();
 FILLCELL_X4 FILLER_72_627 ();
 FILLCELL_X8 FILLER_72_632 ();
 FILLCELL_X4 FILLER_72_640 ();
 FILLCELL_X1 FILLER_72_644 ();
 FILLCELL_X2 FILLER_72_649 ();
 FILLCELL_X2 FILLER_72_737 ();
 FILLCELL_X1 FILLER_72_739 ();
 FILLCELL_X2 FILLER_72_762 ();
 FILLCELL_X2 FILLER_72_789 ();
 FILLCELL_X32 FILLER_72_834 ();
 FILLCELL_X2 FILLER_72_872 ();
 FILLCELL_X1 FILLER_72_874 ();
 FILLCELL_X4 FILLER_72_990 ();
 FILLCELL_X2 FILLER_72_994 ();
 FILLCELL_X1 FILLER_72_1012 ();
 FILLCELL_X8 FILLER_72_1020 ();
 FILLCELL_X2 FILLER_72_1028 ();
 FILLCELL_X1 FILLER_72_1030 ();
 FILLCELL_X4 FILLER_72_1038 ();
 FILLCELL_X2 FILLER_72_1042 ();
 FILLCELL_X2 FILLER_72_1058 ();
 FILLCELL_X1 FILLER_72_1068 ();
 FILLCELL_X1 FILLER_72_1090 ();
 FILLCELL_X1 FILLER_72_1106 ();
 FILLCELL_X4 FILLER_72_1111 ();
 FILLCELL_X1 FILLER_72_1115 ();
 FILLCELL_X4 FILLER_72_1121 ();
 FILLCELL_X1 FILLER_72_1129 ();
 FILLCELL_X8 FILLER_72_1134 ();
 FILLCELL_X1 FILLER_72_1146 ();
 FILLCELL_X8 FILLER_72_1178 ();
 FILLCELL_X4 FILLER_72_1186 ();
 FILLCELL_X2 FILLER_72_1190 ();
 FILLCELL_X1 FILLER_72_1192 ();
 FILLCELL_X8 FILLER_72_1199 ();
 FILLCELL_X2 FILLER_72_1207 ();
 FILLCELL_X32 FILLER_73_1 ();
 FILLCELL_X8 FILLER_73_33 ();
 FILLCELL_X2 FILLER_73_41 ();
 FILLCELL_X8 FILLER_73_62 ();
 FILLCELL_X1 FILLER_73_70 ();
 FILLCELL_X2 FILLER_73_104 ();
 FILLCELL_X2 FILLER_73_129 ();
 FILLCELL_X2 FILLER_73_139 ();
 FILLCELL_X1 FILLER_73_151 ();
 FILLCELL_X1 FILLER_73_159 ();
 FILLCELL_X2 FILLER_73_167 ();
 FILLCELL_X1 FILLER_73_183 ();
 FILLCELL_X8 FILLER_73_187 ();
 FILLCELL_X1 FILLER_73_195 ();
 FILLCELL_X2 FILLER_73_213 ();
 FILLCELL_X1 FILLER_73_215 ();
 FILLCELL_X1 FILLER_73_223 ();
 FILLCELL_X1 FILLER_73_239 ();
 FILLCELL_X4 FILLER_73_253 ();
 FILLCELL_X2 FILLER_73_257 ();
 FILLCELL_X1 FILLER_73_259 ();
 FILLCELL_X16 FILLER_73_273 ();
 FILLCELL_X2 FILLER_73_289 ();
 FILLCELL_X1 FILLER_73_291 ();
 FILLCELL_X1 FILLER_73_325 ();
 FILLCELL_X4 FILLER_73_332 ();
 FILLCELL_X2 FILLER_73_336 ();
 FILLCELL_X4 FILLER_73_345 ();
 FILLCELL_X2 FILLER_73_349 ();
 FILLCELL_X8 FILLER_73_381 ();
 FILLCELL_X4 FILLER_73_389 ();
 FILLCELL_X2 FILLER_73_393 ();
 FILLCELL_X1 FILLER_73_395 ();
 FILLCELL_X1 FILLER_73_403 ();
 FILLCELL_X8 FILLER_73_414 ();
 FILLCELL_X4 FILLER_73_422 ();
 FILLCELL_X8 FILLER_73_430 ();
 FILLCELL_X4 FILLER_73_438 ();
 FILLCELL_X2 FILLER_73_467 ();
 FILLCELL_X1 FILLER_73_481 ();
 FILLCELL_X8 FILLER_73_485 ();
 FILLCELL_X4 FILLER_73_493 ();
 FILLCELL_X8 FILLER_73_510 ();
 FILLCELL_X1 FILLER_73_596 ();
 FILLCELL_X2 FILLER_73_610 ();
 FILLCELL_X1 FILLER_73_612 ();
 FILLCELL_X32 FILLER_73_616 ();
 FILLCELL_X4 FILLER_73_648 ();
 FILLCELL_X8 FILLER_73_655 ();
 FILLCELL_X2 FILLER_73_670 ();
 FILLCELL_X4 FILLER_73_691 ();
 FILLCELL_X8 FILLER_73_699 ();
 FILLCELL_X1 FILLER_73_707 ();
 FILLCELL_X16 FILLER_73_725 ();
 FILLCELL_X2 FILLER_73_741 ();
 FILLCELL_X1 FILLER_73_743 ();
 FILLCELL_X2 FILLER_73_755 ();
 FILLCELL_X1 FILLER_73_757 ();
 FILLCELL_X1 FILLER_73_762 ();
 FILLCELL_X2 FILLER_73_774 ();
 FILLCELL_X1 FILLER_73_811 ();
 FILLCELL_X16 FILLER_73_824 ();
 FILLCELL_X8 FILLER_73_840 ();
 FILLCELL_X4 FILLER_73_960 ();
 FILLCELL_X2 FILLER_73_971 ();
 FILLCELL_X8 FILLER_73_985 ();
 FILLCELL_X2 FILLER_73_993 ();
 FILLCELL_X8 FILLER_73_1019 ();
 FILLCELL_X1 FILLER_73_1027 ();
 FILLCELL_X2 FILLER_73_1044 ();
 FILLCELL_X2 FILLER_73_1051 ();
 FILLCELL_X4 FILLER_73_1072 ();
 FILLCELL_X2 FILLER_73_1076 ();
 FILLCELL_X2 FILLER_73_1092 ();
 FILLCELL_X1 FILLER_73_1101 ();
 FILLCELL_X4 FILLER_73_1113 ();
 FILLCELL_X2 FILLER_73_1117 ();
 FILLCELL_X2 FILLER_73_1123 ();
 FILLCELL_X4 FILLER_73_1129 ();
 FILLCELL_X2 FILLER_73_1133 ();
 FILLCELL_X1 FILLER_73_1151 ();
 FILLCELL_X8 FILLER_73_1181 ();
 FILLCELL_X4 FILLER_73_1189 ();
 FILLCELL_X2 FILLER_73_1193 ();
 FILLCELL_X4 FILLER_73_1198 ();
 FILLCELL_X1 FILLER_73_1202 ();
 FILLCELL_X2 FILLER_73_1206 ();
 FILLCELL_X1 FILLER_73_1208 ();
 FILLCELL_X4 FILLER_74_1 ();
 FILLCELL_X8 FILLER_74_9 ();
 FILLCELL_X4 FILLER_74_17 ();
 FILLCELL_X1 FILLER_74_21 ();
 FILLCELL_X1 FILLER_74_26 ();
 FILLCELL_X32 FILLER_74_30 ();
 FILLCELL_X8 FILLER_74_62 ();
 FILLCELL_X2 FILLER_74_70 ();
 FILLCELL_X1 FILLER_74_72 ();
 FILLCELL_X1 FILLER_74_80 ();
 FILLCELL_X1 FILLER_74_110 ();
 FILLCELL_X1 FILLER_74_121 ();
 FILLCELL_X2 FILLER_74_141 ();
 FILLCELL_X2 FILLER_74_147 ();
 FILLCELL_X2 FILLER_74_164 ();
 FILLCELL_X1 FILLER_74_166 ();
 FILLCELL_X16 FILLER_74_171 ();
 FILLCELL_X8 FILLER_74_187 ();
 FILLCELL_X2 FILLER_74_195 ();
 FILLCELL_X1 FILLER_74_215 ();
 FILLCELL_X2 FILLER_74_247 ();
 FILLCELL_X1 FILLER_74_256 ();
 FILLCELL_X16 FILLER_74_266 ();
 FILLCELL_X4 FILLER_74_282 ();
 FILLCELL_X2 FILLER_74_286 ();
 FILLCELL_X1 FILLER_74_288 ();
 FILLCELL_X16 FILLER_74_296 ();
 FILLCELL_X4 FILLER_74_312 ();
 FILLCELL_X1 FILLER_74_316 ();
 FILLCELL_X2 FILLER_74_328 ();
 FILLCELL_X2 FILLER_74_361 ();
 FILLCELL_X1 FILLER_74_369 ();
 FILLCELL_X8 FILLER_74_381 ();
 FILLCELL_X4 FILLER_74_389 ();
 FILLCELL_X2 FILLER_74_393 ();
 FILLCELL_X1 FILLER_74_395 ();
 FILLCELL_X8 FILLER_74_412 ();
 FILLCELL_X8 FILLER_74_444 ();
 FILLCELL_X4 FILLER_74_452 ();
 FILLCELL_X2 FILLER_74_473 ();
 FILLCELL_X4 FILLER_74_485 ();
 FILLCELL_X2 FILLER_74_489 ();
 FILLCELL_X1 FILLER_74_491 ();
 FILLCELL_X1 FILLER_74_564 ();
 FILLCELL_X2 FILLER_74_572 ();
 FILLCELL_X1 FILLER_74_574 ();
 FILLCELL_X2 FILLER_74_611 ();
 FILLCELL_X1 FILLER_74_613 ();
 FILLCELL_X8 FILLER_74_621 ();
 FILLCELL_X2 FILLER_74_629 ();
 FILLCELL_X8 FILLER_74_632 ();
 FILLCELL_X4 FILLER_74_640 ();
 FILLCELL_X2 FILLER_74_644 ();
 FILLCELL_X1 FILLER_74_646 ();
 FILLCELL_X8 FILLER_74_649 ();
 FILLCELL_X4 FILLER_74_657 ();
 FILLCELL_X2 FILLER_74_661 ();
 FILLCELL_X1 FILLER_74_680 ();
 FILLCELL_X2 FILLER_74_688 ();
 FILLCELL_X1 FILLER_74_690 ();
 FILLCELL_X2 FILLER_74_708 ();
 FILLCELL_X1 FILLER_74_747 ();
 FILLCELL_X2 FILLER_74_755 ();
 FILLCELL_X1 FILLER_74_775 ();
 FILLCELL_X4 FILLER_74_794 ();
 FILLCELL_X8 FILLER_74_820 ();
 FILLCELL_X4 FILLER_74_828 ();
 FILLCELL_X1 FILLER_74_832 ();
 FILLCELL_X2 FILLER_74_860 ();
 FILLCELL_X1 FILLER_74_945 ();
 FILLCELL_X4 FILLER_74_959 ();
 FILLCELL_X2 FILLER_74_963 ();
 FILLCELL_X1 FILLER_74_971 ();
 FILLCELL_X2 FILLER_74_994 ();
 FILLCELL_X1 FILLER_74_996 ();
 FILLCELL_X8 FILLER_74_1023 ();
 FILLCELL_X1 FILLER_74_1031 ();
 FILLCELL_X1 FILLER_74_1072 ();
 FILLCELL_X1 FILLER_74_1078 ();
 FILLCELL_X4 FILLER_74_1082 ();
 FILLCELL_X8 FILLER_74_1108 ();
 FILLCELL_X4 FILLER_74_1116 ();
 FILLCELL_X2 FILLER_74_1120 ();
 FILLCELL_X4 FILLER_74_1128 ();
 FILLCELL_X2 FILLER_74_1132 ();
 FILLCELL_X1 FILLER_74_1140 ();
 FILLCELL_X4 FILLER_74_1146 ();
 FILLCELL_X2 FILLER_74_1150 ();
 FILLCELL_X4 FILLER_74_1159 ();
 FILLCELL_X2 FILLER_74_1170 ();
 FILLCELL_X1 FILLER_74_1172 ();
 FILLCELL_X16 FILLER_74_1193 ();
 FILLCELL_X32 FILLER_75_1 ();
 FILLCELL_X32 FILLER_75_33 ();
 FILLCELL_X4 FILLER_75_65 ();
 FILLCELL_X1 FILLER_75_69 ();
 FILLCELL_X2 FILLER_75_83 ();
 FILLCELL_X1 FILLER_75_85 ();
 FILLCELL_X1 FILLER_75_125 ();
 FILLCELL_X2 FILLER_75_133 ();
 FILLCELL_X2 FILLER_75_140 ();
 FILLCELL_X8 FILLER_75_157 ();
 FILLCELL_X2 FILLER_75_165 ();
 FILLCELL_X1 FILLER_75_167 ();
 FILLCELL_X2 FILLER_75_172 ();
 FILLCELL_X4 FILLER_75_209 ();
 FILLCELL_X2 FILLER_75_213 ();
 FILLCELL_X8 FILLER_75_228 ();
 FILLCELL_X1 FILLER_75_236 ();
 FILLCELL_X4 FILLER_75_239 ();
 FILLCELL_X2 FILLER_75_243 ();
 FILLCELL_X2 FILLER_75_256 ();
 FILLCELL_X16 FILLER_75_268 ();
 FILLCELL_X4 FILLER_75_284 ();
 FILLCELL_X4 FILLER_75_297 ();
 FILLCELL_X2 FILLER_75_301 ();
 FILLCELL_X4 FILLER_75_328 ();
 FILLCELL_X2 FILLER_75_332 ();
 FILLCELL_X4 FILLER_75_340 ();
 FILLCELL_X1 FILLER_75_365 ();
 FILLCELL_X2 FILLER_75_380 ();
 FILLCELL_X2 FILLER_75_399 ();
 FILLCELL_X1 FILLER_75_401 ();
 FILLCELL_X1 FILLER_75_433 ();
 FILLCELL_X2 FILLER_75_450 ();
 FILLCELL_X2 FILLER_75_456 ();
 FILLCELL_X1 FILLER_75_458 ();
 FILLCELL_X2 FILLER_75_466 ();
 FILLCELL_X4 FILLER_75_475 ();
 FILLCELL_X4 FILLER_75_485 ();
 FILLCELL_X2 FILLER_75_489 ();
 FILLCELL_X1 FILLER_75_491 ();
 FILLCELL_X16 FILLER_75_502 ();
 FILLCELL_X4 FILLER_75_518 ();
 FILLCELL_X2 FILLER_75_579 ();
 FILLCELL_X1 FILLER_75_581 ();
 FILLCELL_X2 FILLER_75_599 ();
 FILLCELL_X2 FILLER_75_606 ();
 FILLCELL_X1 FILLER_75_608 ();
 FILLCELL_X8 FILLER_75_629 ();
 FILLCELL_X2 FILLER_75_637 ();
 FILLCELL_X1 FILLER_75_658 ();
 FILLCELL_X2 FILLER_75_663 ();
 FILLCELL_X8 FILLER_75_683 ();
 FILLCELL_X2 FILLER_75_691 ();
 FILLCELL_X1 FILLER_75_693 ();
 FILLCELL_X1 FILLER_75_706 ();
 FILLCELL_X1 FILLER_75_752 ();
 FILLCELL_X4 FILLER_75_766 ();
 FILLCELL_X2 FILLER_75_770 ();
 FILLCELL_X1 FILLER_75_772 ();
 FILLCELL_X2 FILLER_75_781 ();
 FILLCELL_X8 FILLER_75_831 ();
 FILLCELL_X4 FILLER_75_839 ();
 FILLCELL_X2 FILLER_75_843 ();
 FILLCELL_X2 FILLER_75_852 ();
 FILLCELL_X2 FILLER_75_860 ();
 FILLCELL_X1 FILLER_75_867 ();
 FILLCELL_X8 FILLER_75_872 ();
 FILLCELL_X2 FILLER_75_880 ();
 FILLCELL_X1 FILLER_75_882 ();
 FILLCELL_X1 FILLER_75_893 ();
 FILLCELL_X2 FILLER_75_917 ();
 FILLCELL_X8 FILLER_75_956 ();
 FILLCELL_X1 FILLER_75_964 ();
 FILLCELL_X2 FILLER_75_972 ();
 FILLCELL_X1 FILLER_75_974 ();
 FILLCELL_X8 FILLER_75_984 ();
 FILLCELL_X32 FILLER_75_997 ();
 FILLCELL_X2 FILLER_75_1042 ();
 FILLCELL_X8 FILLER_75_1058 ();
 FILLCELL_X2 FILLER_75_1066 ();
 FILLCELL_X1 FILLER_75_1072 ();
 FILLCELL_X4 FILLER_75_1078 ();
 FILLCELL_X4 FILLER_75_1084 ();
 FILLCELL_X2 FILLER_75_1088 ();
 FILLCELL_X8 FILLER_75_1095 ();
 FILLCELL_X4 FILLER_75_1103 ();
 FILLCELL_X1 FILLER_75_1107 ();
 FILLCELL_X2 FILLER_75_1111 ();
 FILLCELL_X1 FILLER_75_1113 ();
 FILLCELL_X1 FILLER_75_1118 ();
 FILLCELL_X8 FILLER_75_1123 ();
 FILLCELL_X4 FILLER_75_1131 ();
 FILLCELL_X1 FILLER_75_1139 ();
 FILLCELL_X2 FILLER_75_1160 ();
 FILLCELL_X1 FILLER_75_1162 ();
 FILLCELL_X8 FILLER_75_1170 ();
 FILLCELL_X2 FILLER_75_1178 ();
 FILLCELL_X1 FILLER_75_1180 ();
 FILLCELL_X16 FILLER_75_1191 ();
 FILLCELL_X2 FILLER_75_1207 ();
 FILLCELL_X4 FILLER_76_1 ();
 FILLCELL_X2 FILLER_76_5 ();
 FILLCELL_X8 FILLER_76_27 ();
 FILLCELL_X1 FILLER_76_35 ();
 FILLCELL_X2 FILLER_76_40 ();
 FILLCELL_X1 FILLER_76_42 ();
 FILLCELL_X8 FILLER_76_51 ();
 FILLCELL_X1 FILLER_76_73 ();
 FILLCELL_X1 FILLER_76_113 ();
 FILLCELL_X2 FILLER_76_121 ();
 FILLCELL_X4 FILLER_76_127 ();
 FILLCELL_X2 FILLER_76_131 ();
 FILLCELL_X1 FILLER_76_133 ();
 FILLCELL_X1 FILLER_76_144 ();
 FILLCELL_X4 FILLER_76_156 ();
 FILLCELL_X2 FILLER_76_160 ();
 FILLCELL_X1 FILLER_76_162 ();
 FILLCELL_X1 FILLER_76_213 ();
 FILLCELL_X4 FILLER_76_229 ();
 FILLCELL_X2 FILLER_76_233 ();
 FILLCELL_X1 FILLER_76_235 ();
 FILLCELL_X4 FILLER_76_245 ();
 FILLCELL_X8 FILLER_76_264 ();
 FILLCELL_X2 FILLER_76_272 ();
 FILLCELL_X32 FILLER_76_279 ();
 FILLCELL_X4 FILLER_76_311 ();
 FILLCELL_X2 FILLER_76_315 ();
 FILLCELL_X4 FILLER_76_330 ();
 FILLCELL_X1 FILLER_76_334 ();
 FILLCELL_X2 FILLER_76_345 ();
 FILLCELL_X2 FILLER_76_358 ();
 FILLCELL_X1 FILLER_76_360 ();
 FILLCELL_X2 FILLER_76_371 ();
 FILLCELL_X2 FILLER_76_379 ();
 FILLCELL_X4 FILLER_76_409 ();
 FILLCELL_X2 FILLER_76_413 ();
 FILLCELL_X2 FILLER_76_444 ();
 FILLCELL_X2 FILLER_76_480 ();
 FILLCELL_X8 FILLER_76_511 ();
 FILLCELL_X1 FILLER_76_519 ();
 FILLCELL_X2 FILLER_76_530 ();
 FILLCELL_X1 FILLER_76_532 ();
 FILLCELL_X2 FILLER_76_545 ();
 FILLCELL_X2 FILLER_76_561 ();
 FILLCELL_X4 FILLER_76_570 ();
 FILLCELL_X1 FILLER_76_574 ();
 FILLCELL_X32 FILLER_76_592 ();
 FILLCELL_X4 FILLER_76_624 ();
 FILLCELL_X2 FILLER_76_628 ();
 FILLCELL_X1 FILLER_76_630 ();
 FILLCELL_X16 FILLER_76_632 ();
 FILLCELL_X4 FILLER_76_648 ();
 FILLCELL_X2 FILLER_76_652 ();
 FILLCELL_X1 FILLER_76_654 ();
 FILLCELL_X4 FILLER_76_662 ();
 FILLCELL_X2 FILLER_76_666 ();
 FILLCELL_X4 FILLER_76_677 ();
 FILLCELL_X1 FILLER_76_692 ();
 FILLCELL_X4 FILLER_76_696 ();
 FILLCELL_X2 FILLER_76_700 ();
 FILLCELL_X1 FILLER_76_702 ();
 FILLCELL_X8 FILLER_76_713 ();
 FILLCELL_X2 FILLER_76_721 ();
 FILLCELL_X4 FILLER_76_736 ();
 FILLCELL_X2 FILLER_76_740 ();
 FILLCELL_X8 FILLER_76_749 ();
 FILLCELL_X2 FILLER_76_757 ();
 FILLCELL_X2 FILLER_76_772 ();
 FILLCELL_X2 FILLER_76_781 ();
 FILLCELL_X2 FILLER_76_804 ();
 FILLCELL_X2 FILLER_76_813 ();
 FILLCELL_X4 FILLER_76_846 ();
 FILLCELL_X1 FILLER_76_850 ();
 FILLCELL_X2 FILLER_76_896 ();
 FILLCELL_X1 FILLER_76_916 ();
 FILLCELL_X4 FILLER_76_953 ();
 FILLCELL_X1 FILLER_76_957 ();
 FILLCELL_X2 FILLER_76_979 ();
 FILLCELL_X16 FILLER_76_987 ();
 FILLCELL_X4 FILLER_76_1003 ();
 FILLCELL_X2 FILLER_76_1007 ();
 FILLCELL_X1 FILLER_76_1009 ();
 FILLCELL_X8 FILLER_76_1017 ();
 FILLCELL_X4 FILLER_76_1025 ();
 FILLCELL_X1 FILLER_76_1029 ();
 FILLCELL_X4 FILLER_76_1039 ();
 FILLCELL_X1 FILLER_76_1043 ();
 FILLCELL_X2 FILLER_76_1076 ();
 FILLCELL_X4 FILLER_76_1090 ();
 FILLCELL_X1 FILLER_76_1094 ();
 FILLCELL_X2 FILLER_76_1100 ();
 FILLCELL_X1 FILLER_76_1102 ();
 FILLCELL_X2 FILLER_76_1106 ();
 FILLCELL_X8 FILLER_76_1134 ();
 FILLCELL_X2 FILLER_76_1152 ();
 FILLCELL_X1 FILLER_76_1154 ();
 FILLCELL_X1 FILLER_76_1205 ();
 FILLCELL_X32 FILLER_77_1 ();
 FILLCELL_X2 FILLER_77_33 ();
 FILLCELL_X4 FILLER_77_39 ();
 FILLCELL_X8 FILLER_77_60 ();
 FILLCELL_X2 FILLER_77_68 ();
 FILLCELL_X1 FILLER_77_70 ();
 FILLCELL_X1 FILLER_77_114 ();
 FILLCELL_X4 FILLER_77_123 ();
 FILLCELL_X4 FILLER_77_131 ();
 FILLCELL_X1 FILLER_77_135 ();
 FILLCELL_X1 FILLER_77_140 ();
 FILLCELL_X4 FILLER_77_145 ();
 FILLCELL_X2 FILLER_77_149 ();
 FILLCELL_X1 FILLER_77_151 ();
 FILLCELL_X1 FILLER_77_179 ();
 FILLCELL_X8 FILLER_77_184 ();
 FILLCELL_X4 FILLER_77_192 ();
 FILLCELL_X2 FILLER_77_196 ();
 FILLCELL_X1 FILLER_77_201 ();
 FILLCELL_X2 FILLER_77_220 ();
 FILLCELL_X8 FILLER_77_244 ();
 FILLCELL_X4 FILLER_77_252 ();
 FILLCELL_X8 FILLER_77_263 ();
 FILLCELL_X4 FILLER_77_271 ();
 FILLCELL_X2 FILLER_77_275 ();
 FILLCELL_X1 FILLER_77_277 ();
 FILLCELL_X4 FILLER_77_295 ();
 FILLCELL_X2 FILLER_77_299 ();
 FILLCELL_X1 FILLER_77_301 ();
 FILLCELL_X1 FILLER_77_341 ();
 FILLCELL_X2 FILLER_77_354 ();
 FILLCELL_X2 FILLER_77_365 ();
 FILLCELL_X2 FILLER_77_385 ();
 FILLCELL_X2 FILLER_77_397 ();
 FILLCELL_X4 FILLER_77_419 ();
 FILLCELL_X1 FILLER_77_459 ();
 FILLCELL_X2 FILLER_77_477 ();
 FILLCELL_X1 FILLER_77_488 ();
 FILLCELL_X1 FILLER_77_501 ();
 FILLCELL_X4 FILLER_77_509 ();
 FILLCELL_X1 FILLER_77_513 ();
 FILLCELL_X2 FILLER_77_539 ();
 FILLCELL_X2 FILLER_77_563 ();
 FILLCELL_X1 FILLER_77_565 ();
 FILLCELL_X32 FILLER_77_583 ();
 FILLCELL_X32 FILLER_77_615 ();
 FILLCELL_X4 FILLER_77_651 ();
 FILLCELL_X2 FILLER_77_655 ();
 FILLCELL_X1 FILLER_77_682 ();
 FILLCELL_X8 FILLER_77_692 ();
 FILLCELL_X2 FILLER_77_700 ();
 FILLCELL_X8 FILLER_77_705 ();
 FILLCELL_X2 FILLER_77_713 ();
 FILLCELL_X4 FILLER_77_719 ();
 FILLCELL_X1 FILLER_77_723 ();
 FILLCELL_X4 FILLER_77_729 ();
 FILLCELL_X2 FILLER_77_733 ();
 FILLCELL_X1 FILLER_77_735 ();
 FILLCELL_X4 FILLER_77_750 ();
 FILLCELL_X1 FILLER_77_754 ();
 FILLCELL_X8 FILLER_77_766 ();
 FILLCELL_X2 FILLER_77_774 ();
 FILLCELL_X2 FILLER_77_810 ();
 FILLCELL_X4 FILLER_77_825 ();
 FILLCELL_X1 FILLER_77_829 ();
 FILLCELL_X2 FILLER_77_855 ();
 FILLCELL_X8 FILLER_77_866 ();
 FILLCELL_X1 FILLER_77_874 ();
 FILLCELL_X8 FILLER_77_882 ();
 FILLCELL_X4 FILLER_77_890 ();
 FILLCELL_X4 FILLER_77_901 ();
 FILLCELL_X1 FILLER_77_905 ();
 FILLCELL_X1 FILLER_77_933 ();
 FILLCELL_X8 FILLER_77_985 ();
 FILLCELL_X2 FILLER_77_993 ();
 FILLCELL_X16 FILLER_77_1012 ();
 FILLCELL_X1 FILLER_77_1028 ();
 FILLCELL_X8 FILLER_77_1034 ();
 FILLCELL_X4 FILLER_77_1042 ();
 FILLCELL_X4 FILLER_77_1053 ();
 FILLCELL_X1 FILLER_77_1057 ();
 FILLCELL_X4 FILLER_77_1064 ();
 FILLCELL_X1 FILLER_77_1068 ();
 FILLCELL_X1 FILLER_77_1080 ();
 FILLCELL_X1 FILLER_77_1094 ();
 FILLCELL_X1 FILLER_77_1105 ();
 FILLCELL_X2 FILLER_77_1110 ();
 FILLCELL_X4 FILLER_77_1116 ();
 FILLCELL_X1 FILLER_77_1120 ();
 FILLCELL_X1 FILLER_77_1131 ();
 FILLCELL_X1 FILLER_77_1141 ();
 FILLCELL_X4 FILLER_77_1148 ();
 FILLCELL_X1 FILLER_77_1152 ();
 FILLCELL_X2 FILLER_77_1177 ();
 FILLCELL_X1 FILLER_77_1179 ();
 FILLCELL_X1 FILLER_77_1184 ();
 FILLCELL_X4 FILLER_77_1199 ();
 FILLCELL_X2 FILLER_77_1206 ();
 FILLCELL_X1 FILLER_77_1208 ();
 FILLCELL_X4 FILLER_78_1 ();
 FILLCELL_X2 FILLER_78_5 ();
 FILLCELL_X1 FILLER_78_7 ();
 FILLCELL_X16 FILLER_78_14 ();
 FILLCELL_X4 FILLER_78_30 ();
 FILLCELL_X2 FILLER_78_34 ();
 FILLCELL_X32 FILLER_78_40 ();
 FILLCELL_X4 FILLER_78_72 ();
 FILLCELL_X2 FILLER_78_76 ();
 FILLCELL_X1 FILLER_78_78 ();
 FILLCELL_X1 FILLER_78_96 ();
 FILLCELL_X2 FILLER_78_103 ();
 FILLCELL_X1 FILLER_78_112 ();
 FILLCELL_X8 FILLER_78_124 ();
 FILLCELL_X4 FILLER_78_132 ();
 FILLCELL_X2 FILLER_78_136 ();
 FILLCELL_X8 FILLER_78_142 ();
 FILLCELL_X4 FILLER_78_158 ();
 FILLCELL_X2 FILLER_78_162 ();
 FILLCELL_X1 FILLER_78_164 ();
 FILLCELL_X4 FILLER_78_168 ();
 FILLCELL_X2 FILLER_78_172 ();
 FILLCELL_X1 FILLER_78_181 ();
 FILLCELL_X1 FILLER_78_197 ();
 FILLCELL_X2 FILLER_78_204 ();
 FILLCELL_X1 FILLER_78_234 ();
 FILLCELL_X32 FILLER_78_254 ();
 FILLCELL_X16 FILLER_78_286 ();
 FILLCELL_X8 FILLER_78_302 ();
 FILLCELL_X2 FILLER_78_310 ();
 FILLCELL_X4 FILLER_78_318 ();
 FILLCELL_X1 FILLER_78_322 ();
 FILLCELL_X2 FILLER_78_333 ();
 FILLCELL_X1 FILLER_78_335 ();
 FILLCELL_X1 FILLER_78_342 ();
 FILLCELL_X16 FILLER_78_349 ();
 FILLCELL_X2 FILLER_78_365 ();
 FILLCELL_X4 FILLER_78_390 ();
 FILLCELL_X1 FILLER_78_400 ();
 FILLCELL_X1 FILLER_78_415 ();
 FILLCELL_X1 FILLER_78_435 ();
 FILLCELL_X1 FILLER_78_446 ();
 FILLCELL_X16 FILLER_78_455 ();
 FILLCELL_X2 FILLER_78_471 ();
 FILLCELL_X2 FILLER_78_495 ();
 FILLCELL_X1 FILLER_78_506 ();
 FILLCELL_X1 FILLER_78_520 ();
 FILLCELL_X4 FILLER_78_534 ();
 FILLCELL_X1 FILLER_78_538 ();
 FILLCELL_X16 FILLER_78_546 ();
 FILLCELL_X2 FILLER_78_562 ();
 FILLCELL_X1 FILLER_78_582 ();
 FILLCELL_X1 FILLER_78_588 ();
 FILLCELL_X16 FILLER_78_613 ();
 FILLCELL_X2 FILLER_78_629 ();
 FILLCELL_X16 FILLER_78_632 ();
 FILLCELL_X4 FILLER_78_648 ();
 FILLCELL_X2 FILLER_78_652 ();
 FILLCELL_X16 FILLER_78_658 ();
 FILLCELL_X4 FILLER_78_674 ();
 FILLCELL_X2 FILLER_78_678 ();
 FILLCELL_X1 FILLER_78_680 ();
 FILLCELL_X4 FILLER_78_700 ();
 FILLCELL_X4 FILLER_78_713 ();
 FILLCELL_X2 FILLER_78_717 ();
 FILLCELL_X8 FILLER_78_730 ();
 FILLCELL_X1 FILLER_78_749 ();
 FILLCELL_X8 FILLER_78_754 ();
 FILLCELL_X1 FILLER_78_762 ();
 FILLCELL_X4 FILLER_78_767 ();
 FILLCELL_X2 FILLER_78_771 ();
 FILLCELL_X1 FILLER_78_796 ();
 FILLCELL_X2 FILLER_78_827 ();
 FILLCELL_X1 FILLER_78_829 ();
 FILLCELL_X1 FILLER_78_833 ();
 FILLCELL_X8 FILLER_78_849 ();
 FILLCELL_X1 FILLER_78_857 ();
 FILLCELL_X2 FILLER_78_875 ();
 FILLCELL_X4 FILLER_78_904 ();
 FILLCELL_X2 FILLER_78_908 ();
 FILLCELL_X2 FILLER_78_926 ();
 FILLCELL_X2 FILLER_78_955 ();
 FILLCELL_X4 FILLER_78_974 ();
 FILLCELL_X2 FILLER_78_978 ();
 FILLCELL_X32 FILLER_78_1002 ();
 FILLCELL_X8 FILLER_78_1034 ();
 FILLCELL_X1 FILLER_78_1042 ();
 FILLCELL_X4 FILLER_78_1047 ();
 FILLCELL_X2 FILLER_78_1062 ();
 FILLCELL_X1 FILLER_78_1064 ();
 FILLCELL_X1 FILLER_78_1081 ();
 FILLCELL_X8 FILLER_78_1087 ();
 FILLCELL_X4 FILLER_78_1095 ();
 FILLCELL_X2 FILLER_78_1099 ();
 FILLCELL_X1 FILLER_78_1101 ();
 FILLCELL_X2 FILLER_78_1109 ();
 FILLCELL_X4 FILLER_78_1117 ();
 FILLCELL_X1 FILLER_78_1121 ();
 FILLCELL_X4 FILLER_78_1135 ();
 FILLCELL_X2 FILLER_78_1139 ();
 FILLCELL_X1 FILLER_78_1141 ();
 FILLCELL_X2 FILLER_78_1147 ();
 FILLCELL_X1 FILLER_78_1161 ();
 FILLCELL_X2 FILLER_78_1169 ();
 FILLCELL_X4 FILLER_78_1176 ();
 FILLCELL_X2 FILLER_78_1180 ();
 FILLCELL_X1 FILLER_78_1182 ();
 FILLCELL_X8 FILLER_78_1186 ();
 FILLCELL_X4 FILLER_78_1194 ();
 FILLCELL_X2 FILLER_78_1198 ();
 FILLCELL_X2 FILLER_78_1206 ();
 FILLCELL_X1 FILLER_78_1208 ();
 FILLCELL_X8 FILLER_79_1 ();
 FILLCELL_X2 FILLER_79_9 ();
 FILLCELL_X1 FILLER_79_11 ();
 FILLCELL_X4 FILLER_79_15 ();
 FILLCELL_X2 FILLER_79_22 ();
 FILLCELL_X1 FILLER_79_24 ();
 FILLCELL_X2 FILLER_79_28 ();
 FILLCELL_X1 FILLER_79_30 ();
 FILLCELL_X4 FILLER_79_34 ();
 FILLCELL_X2 FILLER_79_72 ();
 FILLCELL_X1 FILLER_79_95 ();
 FILLCELL_X2 FILLER_79_100 ();
 FILLCELL_X1 FILLER_79_113 ();
 FILLCELL_X1 FILLER_79_126 ();
 FILLCELL_X2 FILLER_79_130 ();
 FILLCELL_X1 FILLER_79_153 ();
 FILLCELL_X2 FILLER_79_158 ();
 FILLCELL_X4 FILLER_79_179 ();
 FILLCELL_X2 FILLER_79_200 ();
 FILLCELL_X2 FILLER_79_218 ();
 FILLCELL_X1 FILLER_79_220 ();
 FILLCELL_X2 FILLER_79_229 ();
 FILLCELL_X1 FILLER_79_235 ();
 FILLCELL_X2 FILLER_79_240 ();
 FILLCELL_X8 FILLER_79_249 ();
 FILLCELL_X4 FILLER_79_257 ();
 FILLCELL_X2 FILLER_79_261 ();
 FILLCELL_X1 FILLER_79_263 ();
 FILLCELL_X16 FILLER_79_273 ();
 FILLCELL_X2 FILLER_79_289 ();
 FILLCELL_X8 FILLER_79_300 ();
 FILLCELL_X1 FILLER_79_308 ();
 FILLCELL_X4 FILLER_79_315 ();
 FILLCELL_X2 FILLER_79_329 ();
 FILLCELL_X1 FILLER_79_331 ();
 FILLCELL_X8 FILLER_79_354 ();
 FILLCELL_X4 FILLER_79_390 ();
 FILLCELL_X1 FILLER_79_394 ();
 FILLCELL_X2 FILLER_79_411 ();
 FILLCELL_X8 FILLER_79_420 ();
 FILLCELL_X2 FILLER_79_438 ();
 FILLCELL_X1 FILLER_79_447 ();
 FILLCELL_X16 FILLER_79_460 ();
 FILLCELL_X2 FILLER_79_476 ();
 FILLCELL_X1 FILLER_79_478 ();
 FILLCELL_X4 FILLER_79_481 ();
 FILLCELL_X1 FILLER_79_498 ();
 FILLCELL_X1 FILLER_79_512 ();
 FILLCELL_X1 FILLER_79_526 ();
 FILLCELL_X1 FILLER_79_536 ();
 FILLCELL_X1 FILLER_79_541 ();
 FILLCELL_X8 FILLER_79_546 ();
 FILLCELL_X4 FILLER_79_562 ();
 FILLCELL_X2 FILLER_79_566 ();
 FILLCELL_X1 FILLER_79_568 ();
 FILLCELL_X1 FILLER_79_593 ();
 FILLCELL_X8 FILLER_79_600 ();
 FILLCELL_X1 FILLER_79_611 ();
 FILLCELL_X8 FILLER_79_619 ();
 FILLCELL_X4 FILLER_79_627 ();
 FILLCELL_X2 FILLER_79_631 ();
 FILLCELL_X1 FILLER_79_685 ();
 FILLCELL_X2 FILLER_79_697 ();
 FILLCELL_X4 FILLER_79_710 ();
 FILLCELL_X1 FILLER_79_754 ();
 FILLCELL_X8 FILLER_79_823 ();
 FILLCELL_X4 FILLER_79_831 ();
 FILLCELL_X1 FILLER_79_835 ();
 FILLCELL_X2 FILLER_79_840 ();
 FILLCELL_X32 FILLER_79_870 ();
 FILLCELL_X8 FILLER_79_902 ();
 FILLCELL_X2 FILLER_79_910 ();
 FILLCELL_X8 FILLER_79_961 ();
 FILLCELL_X1 FILLER_79_986 ();
 FILLCELL_X8 FILLER_79_992 ();
 FILLCELL_X2 FILLER_79_1000 ();
 FILLCELL_X16 FILLER_79_1010 ();
 FILLCELL_X8 FILLER_79_1026 ();
 FILLCELL_X4 FILLER_79_1034 ();
 FILLCELL_X2 FILLER_79_1038 ();
 FILLCELL_X1 FILLER_79_1040 ();
 FILLCELL_X2 FILLER_79_1048 ();
 FILLCELL_X8 FILLER_79_1053 ();
 FILLCELL_X8 FILLER_79_1086 ();
 FILLCELL_X4 FILLER_79_1094 ();
 FILLCELL_X2 FILLER_79_1098 ();
 FILLCELL_X2 FILLER_79_1107 ();
 FILLCELL_X2 FILLER_79_1120 ();
 FILLCELL_X1 FILLER_79_1126 ();
 FILLCELL_X2 FILLER_79_1133 ();
 FILLCELL_X1 FILLER_79_1144 ();
 FILLCELL_X1 FILLER_79_1149 ();
 FILLCELL_X2 FILLER_79_1174 ();
 FILLCELL_X1 FILLER_79_1176 ();
 FILLCELL_X1 FILLER_79_1181 ();
 FILLCELL_X2 FILLER_79_1189 ();
 FILLCELL_X4 FILLER_79_1204 ();
 FILLCELL_X1 FILLER_79_1208 ();
 FILLCELL_X16 FILLER_80_1 ();
 FILLCELL_X8 FILLER_80_17 ();
 FILLCELL_X4 FILLER_80_25 ();
 FILLCELL_X1 FILLER_80_29 ();
 FILLCELL_X32 FILLER_80_34 ();
 FILLCELL_X16 FILLER_80_66 ();
 FILLCELL_X1 FILLER_80_90 ();
 FILLCELL_X8 FILLER_80_95 ();
 FILLCELL_X1 FILLER_80_103 ();
 FILLCELL_X4 FILLER_80_109 ();
 FILLCELL_X1 FILLER_80_151 ();
 FILLCELL_X1 FILLER_80_166 ();
 FILLCELL_X16 FILLER_80_174 ();
 FILLCELL_X4 FILLER_80_190 ();
 FILLCELL_X2 FILLER_80_194 ();
 FILLCELL_X1 FILLER_80_207 ();
 FILLCELL_X1 FILLER_80_218 ();
 FILLCELL_X8 FILLER_80_229 ();
 FILLCELL_X4 FILLER_80_237 ();
 FILLCELL_X1 FILLER_80_241 ();
 FILLCELL_X8 FILLER_80_254 ();
 FILLCELL_X2 FILLER_80_262 ();
 FILLCELL_X1 FILLER_80_264 ();
 FILLCELL_X16 FILLER_80_282 ();
 FILLCELL_X8 FILLER_80_298 ();
 FILLCELL_X4 FILLER_80_306 ();
 FILLCELL_X2 FILLER_80_310 ();
 FILLCELL_X1 FILLER_80_312 ();
 FILLCELL_X1 FILLER_80_336 ();
 FILLCELL_X1 FILLER_80_347 ();
 FILLCELL_X1 FILLER_80_365 ();
 FILLCELL_X2 FILLER_80_380 ();
 FILLCELL_X1 FILLER_80_382 ();
 FILLCELL_X1 FILLER_80_387 ();
 FILLCELL_X1 FILLER_80_401 ();
 FILLCELL_X8 FILLER_80_413 ();
 FILLCELL_X4 FILLER_80_421 ();
 FILLCELL_X2 FILLER_80_425 ();
 FILLCELL_X1 FILLER_80_427 ();
 FILLCELL_X2 FILLER_80_446 ();
 FILLCELL_X2 FILLER_80_452 ();
 FILLCELL_X1 FILLER_80_454 ();
 FILLCELL_X1 FILLER_80_472 ();
 FILLCELL_X1 FILLER_80_527 ();
 FILLCELL_X2 FILLER_80_531 ();
 FILLCELL_X2 FILLER_80_539 ();
 FILLCELL_X2 FILLER_80_571 ();
 FILLCELL_X1 FILLER_80_573 ();
 FILLCELL_X1 FILLER_80_581 ();
 FILLCELL_X4 FILLER_80_587 ();
 FILLCELL_X1 FILLER_80_591 ();
 FILLCELL_X4 FILLER_80_626 ();
 FILLCELL_X1 FILLER_80_630 ();
 FILLCELL_X16 FILLER_80_632 ();
 FILLCELL_X8 FILLER_80_648 ();
 FILLCELL_X4 FILLER_80_656 ();
 FILLCELL_X2 FILLER_80_660 ();
 FILLCELL_X4 FILLER_80_668 ();
 FILLCELL_X8 FILLER_80_679 ();
 FILLCELL_X1 FILLER_80_687 ();
 FILLCELL_X4 FILLER_80_708 ();
 FILLCELL_X4 FILLER_80_722 ();
 FILLCELL_X4 FILLER_80_733 ();
 FILLCELL_X4 FILLER_80_744 ();
 FILLCELL_X2 FILLER_80_762 ();
 FILLCELL_X1 FILLER_80_764 ();
 FILLCELL_X8 FILLER_80_831 ();
 FILLCELL_X4 FILLER_80_839 ();
 FILLCELL_X2 FILLER_80_843 ();
 FILLCELL_X2 FILLER_80_869 ();
 FILLCELL_X2 FILLER_80_878 ();
 FILLCELL_X2 FILLER_80_886 ();
 FILLCELL_X8 FILLER_80_894 ();
 FILLCELL_X2 FILLER_80_906 ();
 FILLCELL_X1 FILLER_80_908 ();
 FILLCELL_X8 FILLER_80_912 ();
 FILLCELL_X4 FILLER_80_920 ();
 FILLCELL_X1 FILLER_80_924 ();
 FILLCELL_X1 FILLER_80_938 ();
 FILLCELL_X32 FILLER_80_973 ();
 FILLCELL_X8 FILLER_80_1005 ();
 FILLCELL_X2 FILLER_80_1013 ();
 FILLCELL_X2 FILLER_80_1043 ();
 FILLCELL_X2 FILLER_80_1061 ();
 FILLCELL_X4 FILLER_80_1074 ();
 FILLCELL_X4 FILLER_80_1082 ();
 FILLCELL_X16 FILLER_80_1093 ();
 FILLCELL_X4 FILLER_80_1109 ();
 FILLCELL_X4 FILLER_80_1120 ();
 FILLCELL_X1 FILLER_80_1124 ();
 FILLCELL_X2 FILLER_80_1129 ();
 FILLCELL_X4 FILLER_80_1141 ();
 FILLCELL_X1 FILLER_80_1145 ();
 FILLCELL_X4 FILLER_80_1149 ();
 FILLCELL_X2 FILLER_80_1153 ();
 FILLCELL_X1 FILLER_80_1155 ();
 FILLCELL_X1 FILLER_80_1167 ();
 FILLCELL_X2 FILLER_80_1178 ();
 FILLCELL_X1 FILLER_80_1180 ();
 FILLCELL_X1 FILLER_80_1185 ();
 FILLCELL_X16 FILLER_80_1189 ();
 FILLCELL_X4 FILLER_80_1205 ();
 FILLCELL_X4 FILLER_81_1 ();
 FILLCELL_X1 FILLER_81_5 ();
 FILLCELL_X4 FILLER_81_15 ();
 FILLCELL_X2 FILLER_81_29 ();
 FILLCELL_X1 FILLER_81_31 ();
 FILLCELL_X8 FILLER_81_56 ();
 FILLCELL_X4 FILLER_81_64 ();
 FILLCELL_X1 FILLER_81_68 ();
 FILLCELL_X4 FILLER_81_82 ();
 FILLCELL_X2 FILLER_81_108 ();
 FILLCELL_X1 FILLER_81_110 ();
 FILLCELL_X1 FILLER_81_129 ();
 FILLCELL_X2 FILLER_81_136 ();
 FILLCELL_X16 FILLER_81_143 ();
 FILLCELL_X2 FILLER_81_159 ();
 FILLCELL_X1 FILLER_81_161 ();
 FILLCELL_X8 FILLER_81_166 ();
 FILLCELL_X8 FILLER_81_178 ();
 FILLCELL_X8 FILLER_81_191 ();
 FILLCELL_X4 FILLER_81_199 ();
 FILLCELL_X2 FILLER_81_203 ();
 FILLCELL_X2 FILLER_81_213 ();
 FILLCELL_X2 FILLER_81_219 ();
 FILLCELL_X2 FILLER_81_228 ();
 FILLCELL_X8 FILLER_81_233 ();
 FILLCELL_X32 FILLER_81_245 ();
 FILLCELL_X2 FILLER_81_277 ();
 FILLCELL_X1 FILLER_81_279 ();
 FILLCELL_X4 FILLER_81_316 ();
 FILLCELL_X4 FILLER_81_327 ();
 FILLCELL_X2 FILLER_81_353 ();
 FILLCELL_X1 FILLER_81_355 ();
 FILLCELL_X4 FILLER_81_363 ();
 FILLCELL_X2 FILLER_81_367 ();
 FILLCELL_X1 FILLER_81_381 ();
 FILLCELL_X4 FILLER_81_389 ();
 FILLCELL_X2 FILLER_81_393 ();
 FILLCELL_X1 FILLER_81_395 ();
 FILLCELL_X2 FILLER_81_405 ();
 FILLCELL_X4 FILLER_81_418 ();
 FILLCELL_X2 FILLER_81_422 ();
 FILLCELL_X4 FILLER_81_431 ();
 FILLCELL_X2 FILLER_81_444 ();
 FILLCELL_X2 FILLER_81_455 ();
 FILLCELL_X1 FILLER_81_457 ();
 FILLCELL_X4 FILLER_81_461 ();
 FILLCELL_X1 FILLER_81_465 ();
 FILLCELL_X1 FILLER_81_470 ();
 FILLCELL_X4 FILLER_81_495 ();
 FILLCELL_X2 FILLER_81_499 ();
 FILLCELL_X1 FILLER_81_511 ();
 FILLCELL_X1 FILLER_81_521 ();
 FILLCELL_X1 FILLER_81_525 ();
 FILLCELL_X2 FILLER_81_539 ();
 FILLCELL_X1 FILLER_81_541 ();
 FILLCELL_X1 FILLER_81_557 ();
 FILLCELL_X2 FILLER_81_563 ();
 FILLCELL_X1 FILLER_81_565 ();
 FILLCELL_X4 FILLER_81_592 ();
 FILLCELL_X1 FILLER_81_596 ();
 FILLCELL_X2 FILLER_81_607 ();
 FILLCELL_X1 FILLER_81_609 ();
 FILLCELL_X8 FILLER_81_625 ();
 FILLCELL_X4 FILLER_81_633 ();
 FILLCELL_X16 FILLER_81_647 ();
 FILLCELL_X4 FILLER_81_663 ();
 FILLCELL_X1 FILLER_81_667 ();
 FILLCELL_X2 FILLER_81_702 ();
 FILLCELL_X4 FILLER_81_722 ();
 FILLCELL_X2 FILLER_81_726 ();
 FILLCELL_X1 FILLER_81_728 ();
 FILLCELL_X2 FILLER_81_761 ();
 FILLCELL_X1 FILLER_81_763 ();
 FILLCELL_X4 FILLER_81_777 ();
 FILLCELL_X1 FILLER_81_781 ();
 FILLCELL_X2 FILLER_81_789 ();
 FILLCELL_X2 FILLER_81_816 ();
 FILLCELL_X8 FILLER_81_826 ();
 FILLCELL_X2 FILLER_81_834 ();
 FILLCELL_X1 FILLER_81_860 ();
 FILLCELL_X1 FILLER_81_887 ();
 FILLCELL_X4 FILLER_81_922 ();
 FILLCELL_X8 FILLER_81_942 ();
 FILLCELL_X2 FILLER_81_950 ();
 FILLCELL_X1 FILLER_81_952 ();
 FILLCELL_X2 FILLER_81_963 ();
 FILLCELL_X2 FILLER_81_989 ();
 FILLCELL_X32 FILLER_81_996 ();
 FILLCELL_X2 FILLER_81_1028 ();
 FILLCELL_X1 FILLER_81_1044 ();
 FILLCELL_X1 FILLER_81_1063 ();
 FILLCELL_X1 FILLER_81_1075 ();
 FILLCELL_X1 FILLER_81_1079 ();
 FILLCELL_X2 FILLER_81_1091 ();
 FILLCELL_X2 FILLER_81_1102 ();
 FILLCELL_X1 FILLER_81_1108 ();
 FILLCELL_X8 FILLER_81_1120 ();
 FILLCELL_X2 FILLER_81_1128 ();
 FILLCELL_X1 FILLER_81_1130 ();
 FILLCELL_X4 FILLER_81_1134 ();
 FILLCELL_X2 FILLER_81_1138 ();
 FILLCELL_X1 FILLER_81_1186 ();
 FILLCELL_X4 FILLER_81_1193 ();
 FILLCELL_X1 FILLER_81_1197 ();
 FILLCELL_X4 FILLER_81_1201 ();
 FILLCELL_X1 FILLER_81_1205 ();
 FILLCELL_X16 FILLER_82_1 ();
 FILLCELL_X32 FILLER_82_20 ();
 FILLCELL_X16 FILLER_82_52 ();
 FILLCELL_X4 FILLER_82_68 ();
 FILLCELL_X4 FILLER_82_89 ();
 FILLCELL_X2 FILLER_82_93 ();
 FILLCELL_X1 FILLER_82_95 ();
 FILLCELL_X2 FILLER_82_109 ();
 FILLCELL_X4 FILLER_82_140 ();
 FILLCELL_X1 FILLER_82_144 ();
 FILLCELL_X1 FILLER_82_149 ();
 FILLCELL_X4 FILLER_82_157 ();
 FILLCELL_X2 FILLER_82_161 ();
 FILLCELL_X1 FILLER_82_167 ();
 FILLCELL_X16 FILLER_82_176 ();
 FILLCELL_X2 FILLER_82_192 ();
 FILLCELL_X8 FILLER_82_202 ();
 FILLCELL_X4 FILLER_82_210 ();
 FILLCELL_X2 FILLER_82_224 ();
 FILLCELL_X1 FILLER_82_226 ();
 FILLCELL_X4 FILLER_82_234 ();
 FILLCELL_X2 FILLER_82_238 ();
 FILLCELL_X1 FILLER_82_240 ();
 FILLCELL_X32 FILLER_82_245 ();
 FILLCELL_X2 FILLER_82_277 ();
 FILLCELL_X1 FILLER_82_279 ();
 FILLCELL_X1 FILLER_82_302 ();
 FILLCELL_X8 FILLER_82_312 ();
 FILLCELL_X4 FILLER_82_329 ();
 FILLCELL_X4 FILLER_82_372 ();
 FILLCELL_X2 FILLER_82_376 ();
 FILLCELL_X16 FILLER_82_391 ();
 FILLCELL_X16 FILLER_82_412 ();
 FILLCELL_X4 FILLER_82_428 ();
 FILLCELL_X2 FILLER_82_451 ();
 FILLCELL_X1 FILLER_82_466 ();
 FILLCELL_X2 FILLER_82_477 ();
 FILLCELL_X4 FILLER_82_488 ();
 FILLCELL_X16 FILLER_82_499 ();
 FILLCELL_X4 FILLER_82_515 ();
 FILLCELL_X1 FILLER_82_519 ();
 FILLCELL_X16 FILLER_82_529 ();
 FILLCELL_X4 FILLER_82_545 ();
 FILLCELL_X1 FILLER_82_549 ();
 FILLCELL_X4 FILLER_82_567 ();
 FILLCELL_X1 FILLER_82_571 ();
 FILLCELL_X8 FILLER_82_582 ();
 FILLCELL_X8 FILLER_82_616 ();
 FILLCELL_X4 FILLER_82_624 ();
 FILLCELL_X2 FILLER_82_628 ();
 FILLCELL_X1 FILLER_82_630 ();
 FILLCELL_X32 FILLER_82_632 ();
 FILLCELL_X8 FILLER_82_664 ();
 FILLCELL_X1 FILLER_82_672 ();
 FILLCELL_X2 FILLER_82_699 ();
 FILLCELL_X4 FILLER_82_708 ();
 FILLCELL_X2 FILLER_82_712 ();
 FILLCELL_X2 FILLER_82_741 ();
 FILLCELL_X4 FILLER_82_750 ();
 FILLCELL_X2 FILLER_82_754 ();
 FILLCELL_X8 FILLER_82_774 ();
 FILLCELL_X1 FILLER_82_782 ();
 FILLCELL_X16 FILLER_82_851 ();
 FILLCELL_X2 FILLER_82_867 ();
 FILLCELL_X8 FILLER_82_895 ();
 FILLCELL_X2 FILLER_82_903 ();
 FILLCELL_X1 FILLER_82_905 ();
 FILLCELL_X2 FILLER_82_912 ();
 FILLCELL_X1 FILLER_82_914 ();
 FILLCELL_X2 FILLER_82_918 ();
 FILLCELL_X4 FILLER_82_937 ();
 FILLCELL_X2 FILLER_82_965 ();
 FILLCELL_X32 FILLER_82_980 ();
 FILLCELL_X16 FILLER_82_1012 ();
 FILLCELL_X8 FILLER_82_1028 ();
 FILLCELL_X2 FILLER_82_1036 ();
 FILLCELL_X2 FILLER_82_1042 ();
 FILLCELL_X1 FILLER_82_1044 ();
 FILLCELL_X1 FILLER_82_1048 ();
 FILLCELL_X4 FILLER_82_1085 ();
 FILLCELL_X2 FILLER_82_1089 ();
 FILLCELL_X8 FILLER_82_1101 ();
 FILLCELL_X1 FILLER_82_1109 ();
 FILLCELL_X4 FILLER_82_1117 ();
 FILLCELL_X2 FILLER_82_1139 ();
 FILLCELL_X1 FILLER_82_1141 ();
 FILLCELL_X8 FILLER_82_1150 ();
 FILLCELL_X1 FILLER_82_1158 ();
 FILLCELL_X2 FILLER_82_1170 ();
 FILLCELL_X1 FILLER_82_1172 ();
 FILLCELL_X1 FILLER_82_1177 ();
 FILLCELL_X2 FILLER_82_1182 ();
 FILLCELL_X8 FILLER_82_1197 ();
 FILLCELL_X4 FILLER_82_1205 ();
 FILLCELL_X4 FILLER_83_1 ();
 FILLCELL_X2 FILLER_83_5 ();
 FILLCELL_X1 FILLER_83_7 ();
 FILLCELL_X8 FILLER_83_12 ();
 FILLCELL_X4 FILLER_83_20 ();
 FILLCELL_X16 FILLER_83_52 ();
 FILLCELL_X8 FILLER_83_85 ();
 FILLCELL_X2 FILLER_83_101 ();
 FILLCELL_X2 FILLER_83_111 ();
 FILLCELL_X1 FILLER_83_113 ();
 FILLCELL_X1 FILLER_83_131 ();
 FILLCELL_X2 FILLER_83_148 ();
 FILLCELL_X1 FILLER_83_150 ();
 FILLCELL_X4 FILLER_83_162 ();
 FILLCELL_X1 FILLER_83_171 ();
 FILLCELL_X8 FILLER_83_175 ();
 FILLCELL_X1 FILLER_83_183 ();
 FILLCELL_X4 FILLER_83_199 ();
 FILLCELL_X1 FILLER_83_206 ();
 FILLCELL_X4 FILLER_83_211 ();
 FILLCELL_X2 FILLER_83_215 ();
 FILLCELL_X8 FILLER_83_232 ();
 FILLCELL_X2 FILLER_83_240 ();
 FILLCELL_X8 FILLER_83_249 ();
 FILLCELL_X4 FILLER_83_257 ();
 FILLCELL_X2 FILLER_83_261 ();
 FILLCELL_X1 FILLER_83_263 ();
 FILLCELL_X8 FILLER_83_273 ();
 FILLCELL_X2 FILLER_83_291 ();
 FILLCELL_X1 FILLER_83_293 ();
 FILLCELL_X2 FILLER_83_335 ();
 FILLCELL_X4 FILLER_83_343 ();
 FILLCELL_X1 FILLER_83_351 ();
 FILLCELL_X2 FILLER_83_354 ();
 FILLCELL_X4 FILLER_83_378 ();
 FILLCELL_X2 FILLER_83_382 ();
 FILLCELL_X1 FILLER_83_384 ();
 FILLCELL_X8 FILLER_83_392 ();
 FILLCELL_X1 FILLER_83_417 ();
 FILLCELL_X4 FILLER_83_421 ();
 FILLCELL_X2 FILLER_83_425 ();
 FILLCELL_X2 FILLER_83_475 ();
 FILLCELL_X1 FILLER_83_494 ();
 FILLCELL_X4 FILLER_83_514 ();
 FILLCELL_X2 FILLER_83_518 ();
 FILLCELL_X4 FILLER_83_536 ();
 FILLCELL_X2 FILLER_83_540 ();
 FILLCELL_X4 FILLER_83_559 ();
 FILLCELL_X2 FILLER_83_570 ();
 FILLCELL_X1 FILLER_83_572 ();
 FILLCELL_X1 FILLER_83_582 ();
 FILLCELL_X16 FILLER_83_585 ();
 FILLCELL_X1 FILLER_83_601 ();
 FILLCELL_X8 FILLER_83_630 ();
 FILLCELL_X4 FILLER_83_638 ();
 FILLCELL_X2 FILLER_83_642 ();
 FILLCELL_X1 FILLER_83_644 ();
 FILLCELL_X8 FILLER_83_652 ();
 FILLCELL_X4 FILLER_83_660 ();
 FILLCELL_X2 FILLER_83_664 ();
 FILLCELL_X32 FILLER_83_690 ();
 FILLCELL_X8 FILLER_83_722 ();
 FILLCELL_X4 FILLER_83_730 ();
 FILLCELL_X2 FILLER_83_734 ();
 FILLCELL_X8 FILLER_83_767 ();
 FILLCELL_X4 FILLER_83_775 ();
 FILLCELL_X2 FILLER_83_779 ();
 FILLCELL_X2 FILLER_83_833 ();
 FILLCELL_X1 FILLER_83_835 ();
 FILLCELL_X4 FILLER_83_860 ();
 FILLCELL_X2 FILLER_83_864 ();
 FILLCELL_X4 FILLER_83_900 ();
 FILLCELL_X1 FILLER_83_904 ();
 FILLCELL_X2 FILLER_83_928 ();
 FILLCELL_X1 FILLER_83_937 ();
 FILLCELL_X1 FILLER_83_944 ();
 FILLCELL_X16 FILLER_83_955 ();
 FILLCELL_X1 FILLER_83_971 ();
 FILLCELL_X1 FILLER_83_978 ();
 FILLCELL_X4 FILLER_83_1000 ();
 FILLCELL_X1 FILLER_83_1004 ();
 FILLCELL_X16 FILLER_83_1014 ();
 FILLCELL_X4 FILLER_83_1030 ();
 FILLCELL_X2 FILLER_83_1034 ();
 FILLCELL_X1 FILLER_83_1036 ();
 FILLCELL_X2 FILLER_83_1059 ();
 FILLCELL_X1 FILLER_83_1061 ();
 FILLCELL_X1 FILLER_83_1075 ();
 FILLCELL_X2 FILLER_83_1080 ();
 FILLCELL_X1 FILLER_83_1082 ();
 FILLCELL_X1 FILLER_83_1086 ();
 FILLCELL_X2 FILLER_83_1091 ();
 FILLCELL_X1 FILLER_83_1093 ();
 FILLCELL_X2 FILLER_83_1098 ();
 FILLCELL_X1 FILLER_83_1100 ();
 FILLCELL_X8 FILLER_83_1105 ();
 FILLCELL_X4 FILLER_83_1113 ();
 FILLCELL_X4 FILLER_83_1132 ();
 FILLCELL_X2 FILLER_83_1136 ();
 FILLCELL_X4 FILLER_83_1161 ();
 FILLCELL_X1 FILLER_83_1165 ();
 FILLCELL_X2 FILLER_83_1171 ();
 FILLCELL_X1 FILLER_83_1187 ();
 FILLCELL_X8 FILLER_83_1191 ();
 FILLCELL_X2 FILLER_83_1199 ();
 FILLCELL_X2 FILLER_83_1204 ();
 FILLCELL_X16 FILLER_84_1 ();
 FILLCELL_X4 FILLER_84_17 ();
 FILLCELL_X1 FILLER_84_21 ();
 FILLCELL_X32 FILLER_84_25 ();
 FILLCELL_X1 FILLER_84_57 ();
 FILLCELL_X8 FILLER_84_66 ();
 FILLCELL_X4 FILLER_84_74 ();
 FILLCELL_X2 FILLER_84_78 ();
 FILLCELL_X2 FILLER_84_100 ();
 FILLCELL_X4 FILLER_84_111 ();
 FILLCELL_X2 FILLER_84_115 ();
 FILLCELL_X2 FILLER_84_121 ();
 FILLCELL_X1 FILLER_84_123 ();
 FILLCELL_X8 FILLER_84_128 ();
 FILLCELL_X16 FILLER_84_141 ();
 FILLCELL_X1 FILLER_84_157 ();
 FILLCELL_X1 FILLER_84_169 ();
 FILLCELL_X1 FILLER_84_177 ();
 FILLCELL_X2 FILLER_84_182 ();
 FILLCELL_X1 FILLER_84_184 ();
 FILLCELL_X8 FILLER_84_191 ();
 FILLCELL_X4 FILLER_84_199 ();
 FILLCELL_X1 FILLER_84_211 ();
 FILLCELL_X1 FILLER_84_222 ();
 FILLCELL_X1 FILLER_84_228 ();
 FILLCELL_X4 FILLER_84_233 ();
 FILLCELL_X32 FILLER_84_243 ();
 FILLCELL_X8 FILLER_84_275 ();
 FILLCELL_X4 FILLER_84_283 ();
 FILLCELL_X2 FILLER_84_287 ();
 FILLCELL_X2 FILLER_84_324 ();
 FILLCELL_X1 FILLER_84_326 ();
 FILLCELL_X8 FILLER_84_337 ();
 FILLCELL_X1 FILLER_84_349 ();
 FILLCELL_X2 FILLER_84_370 ();
 FILLCELL_X1 FILLER_84_372 ();
 FILLCELL_X2 FILLER_84_396 ();
 FILLCELL_X2 FILLER_84_405 ();
 FILLCELL_X1 FILLER_84_416 ();
 FILLCELL_X1 FILLER_84_420 ();
 FILLCELL_X2 FILLER_84_452 ();
 FILLCELL_X1 FILLER_84_454 ();
 FILLCELL_X4 FILLER_84_484 ();
 FILLCELL_X1 FILLER_84_488 ();
 FILLCELL_X2 FILLER_84_501 ();
 FILLCELL_X8 FILLER_84_509 ();
 FILLCELL_X2 FILLER_84_517 ();
 FILLCELL_X1 FILLER_84_519 ();
 FILLCELL_X8 FILLER_84_564 ();
 FILLCELL_X2 FILLER_84_572 ();
 FILLCELL_X1 FILLER_84_574 ();
 FILLCELL_X1 FILLER_84_580 ();
 FILLCELL_X2 FILLER_84_590 ();
 FILLCELL_X4 FILLER_84_595 ();
 FILLCELL_X2 FILLER_84_599 ();
 FILLCELL_X4 FILLER_84_625 ();
 FILLCELL_X2 FILLER_84_629 ();
 FILLCELL_X2 FILLER_84_632 ();
 FILLCELL_X8 FILLER_84_663 ();
 FILLCELL_X4 FILLER_84_671 ();
 FILLCELL_X8 FILLER_84_684 ();
 FILLCELL_X4 FILLER_84_706 ();
 FILLCELL_X1 FILLER_84_710 ();
 FILLCELL_X1 FILLER_84_733 ();
 FILLCELL_X8 FILLER_84_747 ();
 FILLCELL_X4 FILLER_84_755 ();
 FILLCELL_X2 FILLER_84_759 ();
 FILLCELL_X16 FILLER_84_774 ();
 FILLCELL_X1 FILLER_84_790 ();
 FILLCELL_X2 FILLER_84_795 ();
 FILLCELL_X1 FILLER_84_800 ();
 FILLCELL_X8 FILLER_84_805 ();
 FILLCELL_X4 FILLER_84_813 ();
 FILLCELL_X1 FILLER_84_817 ();
 FILLCELL_X1 FILLER_84_832 ();
 FILLCELL_X1 FILLER_84_882 ();
 FILLCELL_X8 FILLER_84_906 ();
 FILLCELL_X8 FILLER_84_957 ();
 FILLCELL_X4 FILLER_84_965 ();
 FILLCELL_X2 FILLER_84_969 ();
 FILLCELL_X16 FILLER_84_981 ();
 FILLCELL_X4 FILLER_84_997 ();
 FILLCELL_X2 FILLER_84_1001 ();
 FILLCELL_X2 FILLER_84_1044 ();
 FILLCELL_X1 FILLER_84_1046 ();
 FILLCELL_X4 FILLER_84_1062 ();
 FILLCELL_X1 FILLER_84_1070 ();
 FILLCELL_X1 FILLER_84_1075 ();
 FILLCELL_X2 FILLER_84_1080 ();
 FILLCELL_X1 FILLER_84_1082 ();
 FILLCELL_X4 FILLER_84_1098 ();
 FILLCELL_X2 FILLER_84_1106 ();
 FILLCELL_X1 FILLER_84_1108 ();
 FILLCELL_X4 FILLER_84_1113 ();
 FILLCELL_X4 FILLER_84_1120 ();
 FILLCELL_X2 FILLER_84_1124 ();
 FILLCELL_X8 FILLER_84_1129 ();
 FILLCELL_X2 FILLER_84_1137 ();
 FILLCELL_X4 FILLER_84_1149 ();
 FILLCELL_X2 FILLER_84_1153 ();
 FILLCELL_X1 FILLER_84_1155 ();
 FILLCELL_X8 FILLER_84_1183 ();
 FILLCELL_X2 FILLER_84_1191 ();
 FILLCELL_X8 FILLER_84_1197 ();
 FILLCELL_X4 FILLER_84_1205 ();
 FILLCELL_X16 FILLER_85_1 ();
 FILLCELL_X8 FILLER_85_17 ();
 FILLCELL_X2 FILLER_85_25 ();
 FILLCELL_X1 FILLER_85_27 ();
 FILLCELL_X16 FILLER_85_35 ();
 FILLCELL_X4 FILLER_85_51 ();
 FILLCELL_X2 FILLER_85_55 ();
 FILLCELL_X8 FILLER_85_74 ();
 FILLCELL_X2 FILLER_85_82 ();
 FILLCELL_X1 FILLER_85_84 ();
 FILLCELL_X2 FILLER_85_105 ();
 FILLCELL_X1 FILLER_85_107 ();
 FILLCELL_X1 FILLER_85_112 ();
 FILLCELL_X1 FILLER_85_123 ();
 FILLCELL_X8 FILLER_85_152 ();
 FILLCELL_X4 FILLER_85_160 ();
 FILLCELL_X2 FILLER_85_164 ();
 FILLCELL_X2 FILLER_85_173 ();
 FILLCELL_X1 FILLER_85_175 ();
 FILLCELL_X2 FILLER_85_179 ();
 FILLCELL_X4 FILLER_85_186 ();
 FILLCELL_X1 FILLER_85_190 ();
 FILLCELL_X4 FILLER_85_206 ();
 FILLCELL_X2 FILLER_85_219 ();
 FILLCELL_X1 FILLER_85_236 ();
 FILLCELL_X8 FILLER_85_246 ();
 FILLCELL_X2 FILLER_85_254 ();
 FILLCELL_X1 FILLER_85_256 ();
 FILLCELL_X16 FILLER_85_276 ();
 FILLCELL_X2 FILLER_85_292 ();
 FILLCELL_X1 FILLER_85_294 ();
 FILLCELL_X4 FILLER_85_320 ();
 FILLCELL_X1 FILLER_85_324 ();
 FILLCELL_X4 FILLER_85_340 ();
 FILLCELL_X8 FILLER_85_352 ();
 FILLCELL_X2 FILLER_85_360 ();
 FILLCELL_X2 FILLER_85_391 ();
 FILLCELL_X2 FILLER_85_407 ();
 FILLCELL_X2 FILLER_85_416 ();
 FILLCELL_X2 FILLER_85_445 ();
 FILLCELL_X4 FILLER_85_478 ();
 FILLCELL_X2 FILLER_85_482 ();
 FILLCELL_X1 FILLER_85_484 ();
 FILLCELL_X4 FILLER_85_488 ();
 FILLCELL_X4 FILLER_85_541 ();
 FILLCELL_X2 FILLER_85_545 ();
 FILLCELL_X8 FILLER_85_563 ();
 FILLCELL_X1 FILLER_85_571 ();
 FILLCELL_X8 FILLER_85_603 ();
 FILLCELL_X1 FILLER_85_611 ();
 FILLCELL_X8 FILLER_85_622 ();
 FILLCELL_X2 FILLER_85_630 ();
 FILLCELL_X8 FILLER_85_639 ();
 FILLCELL_X1 FILLER_85_647 ();
 FILLCELL_X4 FILLER_85_666 ();
 FILLCELL_X1 FILLER_85_670 ();
 FILLCELL_X16 FILLER_85_676 ();
 FILLCELL_X1 FILLER_85_692 ();
 FILLCELL_X16 FILLER_85_704 ();
 FILLCELL_X1 FILLER_85_720 ();
 FILLCELL_X1 FILLER_85_728 ();
 FILLCELL_X4 FILLER_85_758 ();
 FILLCELL_X2 FILLER_85_762 ();
 FILLCELL_X8 FILLER_85_767 ();
 FILLCELL_X4 FILLER_85_775 ();
 FILLCELL_X4 FILLER_85_814 ();
 FILLCELL_X4 FILLER_85_845 ();
 FILLCELL_X2 FILLER_85_849 ();
 FILLCELL_X1 FILLER_85_851 ();
 FILLCELL_X1 FILLER_85_861 ();
 FILLCELL_X4 FILLER_85_916 ();
 FILLCELL_X2 FILLER_85_930 ();
 FILLCELL_X4 FILLER_85_942 ();
 FILLCELL_X2 FILLER_85_946 ();
 FILLCELL_X32 FILLER_85_972 ();
 FILLCELL_X16 FILLER_85_1004 ();
 FILLCELL_X2 FILLER_85_1020 ();
 FILLCELL_X1 FILLER_85_1022 ();
 FILLCELL_X4 FILLER_85_1029 ();
 FILLCELL_X1 FILLER_85_1033 ();
 FILLCELL_X4 FILLER_85_1048 ();
 FILLCELL_X2 FILLER_85_1052 ();
 FILLCELL_X2 FILLER_85_1070 ();
 FILLCELL_X2 FILLER_85_1090 ();
 FILLCELL_X2 FILLER_85_1098 ();
 FILLCELL_X8 FILLER_85_1103 ();
 FILLCELL_X1 FILLER_85_1114 ();
 FILLCELL_X4 FILLER_85_1119 ();
 FILLCELL_X2 FILLER_85_1127 ();
 FILLCELL_X1 FILLER_85_1129 ();
 FILLCELL_X4 FILLER_85_1134 ();
 FILLCELL_X1 FILLER_85_1138 ();
 FILLCELL_X1 FILLER_85_1169 ();
 FILLCELL_X1 FILLER_85_1187 ();
 FILLCELL_X4 FILLER_85_1191 ();
 FILLCELL_X2 FILLER_85_1195 ();
 FILLCELL_X2 FILLER_85_1200 ();
 FILLCELL_X1 FILLER_85_1202 ();
 FILLCELL_X2 FILLER_85_1207 ();
 FILLCELL_X8 FILLER_86_1 ();
 FILLCELL_X2 FILLER_86_9 ();
 FILLCELL_X8 FILLER_86_14 ();
 FILLCELL_X32 FILLER_86_26 ();
 FILLCELL_X16 FILLER_86_58 ();
 FILLCELL_X8 FILLER_86_74 ();
 FILLCELL_X4 FILLER_86_82 ();
 FILLCELL_X1 FILLER_86_86 ();
 FILLCELL_X2 FILLER_86_100 ();
 FILLCELL_X1 FILLER_86_102 ();
 FILLCELL_X1 FILLER_86_107 ();
 FILLCELL_X2 FILLER_86_118 ();
 FILLCELL_X1 FILLER_86_120 ();
 FILLCELL_X4 FILLER_86_124 ();
 FILLCELL_X2 FILLER_86_136 ();
 FILLCELL_X1 FILLER_86_138 ();
 FILLCELL_X8 FILLER_86_145 ();
 FILLCELL_X2 FILLER_86_161 ();
 FILLCELL_X1 FILLER_86_163 ();
 FILLCELL_X4 FILLER_86_175 ();
 FILLCELL_X8 FILLER_86_183 ();
 FILLCELL_X2 FILLER_86_191 ();
 FILLCELL_X16 FILLER_86_197 ();
 FILLCELL_X2 FILLER_86_213 ();
 FILLCELL_X1 FILLER_86_215 ();
 FILLCELL_X1 FILLER_86_220 ();
 FILLCELL_X1 FILLER_86_225 ();
 FILLCELL_X1 FILLER_86_230 ();
 FILLCELL_X1 FILLER_86_238 ();
 FILLCELL_X32 FILLER_86_245 ();
 FILLCELL_X16 FILLER_86_277 ();
 FILLCELL_X8 FILLER_86_293 ();
 FILLCELL_X4 FILLER_86_301 ();
 FILLCELL_X1 FILLER_86_305 ();
 FILLCELL_X1 FILLER_86_312 ();
 FILLCELL_X1 FILLER_86_319 ();
 FILLCELL_X1 FILLER_86_326 ();
 FILLCELL_X8 FILLER_86_333 ();
 FILLCELL_X2 FILLER_86_341 ();
 FILLCELL_X1 FILLER_86_343 ();
 FILLCELL_X2 FILLER_86_357 ();
 FILLCELL_X1 FILLER_86_372 ();
 FILLCELL_X1 FILLER_86_379 ();
 FILLCELL_X8 FILLER_86_406 ();
 FILLCELL_X4 FILLER_86_414 ();
 FILLCELL_X2 FILLER_86_452 ();
 FILLCELL_X8 FILLER_86_476 ();
 FILLCELL_X4 FILLER_86_484 ();
 FILLCELL_X2 FILLER_86_488 ();
 FILLCELL_X16 FILLER_86_495 ();
 FILLCELL_X8 FILLER_86_511 ();
 FILLCELL_X1 FILLER_86_519 ();
 FILLCELL_X16 FILLER_86_555 ();
 FILLCELL_X8 FILLER_86_571 ();
 FILLCELL_X1 FILLER_86_579 ();
 FILLCELL_X4 FILLER_86_593 ();
 FILLCELL_X1 FILLER_86_597 ();
 FILLCELL_X8 FILLER_86_620 ();
 FILLCELL_X2 FILLER_86_628 ();
 FILLCELL_X1 FILLER_86_630 ();
 FILLCELL_X2 FILLER_86_632 ();
 FILLCELL_X1 FILLER_86_634 ();
 FILLCELL_X8 FILLER_86_644 ();
 FILLCELL_X4 FILLER_86_652 ();
 FILLCELL_X4 FILLER_86_682 ();
 FILLCELL_X2 FILLER_86_695 ();
 FILLCELL_X2 FILLER_86_720 ();
 FILLCELL_X1 FILLER_86_722 ();
 FILLCELL_X8 FILLER_86_732 ();
 FILLCELL_X1 FILLER_86_743 ();
 FILLCELL_X1 FILLER_86_751 ();
 FILLCELL_X4 FILLER_86_759 ();
 FILLCELL_X2 FILLER_86_763 ();
 FILLCELL_X1 FILLER_86_819 ();
 FILLCELL_X1 FILLER_86_837 ();
 FILLCELL_X2 FILLER_86_841 ();
 FILLCELL_X4 FILLER_86_854 ();
 FILLCELL_X1 FILLER_86_871 ();
 FILLCELL_X2 FILLER_86_893 ();
 FILLCELL_X4 FILLER_86_929 ();
 FILLCELL_X1 FILLER_86_949 ();
 FILLCELL_X1 FILLER_86_956 ();
 FILLCELL_X2 FILLER_86_976 ();
 FILLCELL_X16 FILLER_86_984 ();
 FILLCELL_X4 FILLER_86_1000 ();
 FILLCELL_X2 FILLER_86_1004 ();
 FILLCELL_X16 FILLER_86_1023 ();
 FILLCELL_X8 FILLER_86_1039 ();
 FILLCELL_X2 FILLER_86_1047 ();
 FILLCELL_X1 FILLER_86_1072 ();
 FILLCELL_X1 FILLER_86_1078 ();
 FILLCELL_X4 FILLER_86_1103 ();
 FILLCELL_X2 FILLER_86_1107 ();
 FILLCELL_X1 FILLER_86_1109 ();
 FILLCELL_X1 FILLER_86_1143 ();
 FILLCELL_X2 FILLER_86_1148 ();
 FILLCELL_X1 FILLER_86_1150 ();
 FILLCELL_X2 FILLER_86_1162 ();
 FILLCELL_X1 FILLER_86_1164 ();
 FILLCELL_X2 FILLER_86_1181 ();
 FILLCELL_X1 FILLER_86_1183 ();
 FILLCELL_X8 FILLER_86_1187 ();
 FILLCELL_X2 FILLER_86_1195 ();
 FILLCELL_X4 FILLER_86_1204 ();
 FILLCELL_X1 FILLER_86_1208 ();
 FILLCELL_X16 FILLER_87_1 ();
 FILLCELL_X1 FILLER_87_17 ();
 FILLCELL_X4 FILLER_87_24 ();
 FILLCELL_X2 FILLER_87_28 ();
 FILLCELL_X32 FILLER_87_33 ();
 FILLCELL_X16 FILLER_87_65 ();
 FILLCELL_X8 FILLER_87_108 ();
 FILLCELL_X2 FILLER_87_116 ();
 FILLCELL_X2 FILLER_87_133 ();
 FILLCELL_X16 FILLER_87_143 ();
 FILLCELL_X8 FILLER_87_159 ();
 FILLCELL_X4 FILLER_87_167 ();
 FILLCELL_X4 FILLER_87_182 ();
 FILLCELL_X2 FILLER_87_186 ();
 FILLCELL_X2 FILLER_87_213 ();
 FILLCELL_X1 FILLER_87_215 ();
 FILLCELL_X1 FILLER_87_221 ();
 FILLCELL_X1 FILLER_87_226 ();
 FILLCELL_X2 FILLER_87_235 ();
 FILLCELL_X1 FILLER_87_237 ();
 FILLCELL_X1 FILLER_87_241 ();
 FILLCELL_X16 FILLER_87_251 ();
 FILLCELL_X8 FILLER_87_267 ();
 FILLCELL_X2 FILLER_87_275 ();
 FILLCELL_X16 FILLER_87_286 ();
 FILLCELL_X1 FILLER_87_308 ();
 FILLCELL_X1 FILLER_87_315 ();
 FILLCELL_X4 FILLER_87_322 ();
 FILLCELL_X2 FILLER_87_326 ();
 FILLCELL_X1 FILLER_87_328 ();
 FILLCELL_X2 FILLER_87_345 ();
 FILLCELL_X1 FILLER_87_347 ();
 FILLCELL_X2 FILLER_87_368 ();
 FILLCELL_X1 FILLER_87_376 ();
 FILLCELL_X4 FILLER_87_405 ();
 FILLCELL_X1 FILLER_87_409 ();
 FILLCELL_X4 FILLER_87_416 ();
 FILLCELL_X2 FILLER_87_420 ();
 FILLCELL_X1 FILLER_87_432 ();
 FILLCELL_X8 FILLER_87_456 ();
 FILLCELL_X32 FILLER_87_542 ();
 FILLCELL_X4 FILLER_87_574 ();
 FILLCELL_X1 FILLER_87_578 ();
 FILLCELL_X2 FILLER_87_581 ();
 FILLCELL_X4 FILLER_87_605 ();
 FILLCELL_X8 FILLER_87_618 ();
 FILLCELL_X4 FILLER_87_626 ();
 FILLCELL_X2 FILLER_87_630 ();
 FILLCELL_X1 FILLER_87_632 ();
 FILLCELL_X8 FILLER_87_643 ();
 FILLCELL_X2 FILLER_87_651 ();
 FILLCELL_X1 FILLER_87_657 ();
 FILLCELL_X4 FILLER_87_663 ();
 FILLCELL_X1 FILLER_87_667 ();
 FILLCELL_X2 FILLER_87_687 ();
 FILLCELL_X4 FILLER_87_708 ();
 FILLCELL_X4 FILLER_87_721 ();
 FILLCELL_X1 FILLER_87_725 ();
 FILLCELL_X8 FILLER_87_733 ();
 FILLCELL_X2 FILLER_87_741 ();
 FILLCELL_X1 FILLER_87_743 ();
 FILLCELL_X16 FILLER_87_761 ();
 FILLCELL_X1 FILLER_87_777 ();
 FILLCELL_X4 FILLER_87_788 ();
 FILLCELL_X2 FILLER_87_792 ();
 FILLCELL_X1 FILLER_87_794 ();
 FILLCELL_X4 FILLER_87_857 ();
 FILLCELL_X8 FILLER_87_870 ();
 FILLCELL_X2 FILLER_87_900 ();
 FILLCELL_X2 FILLER_87_918 ();
 FILLCELL_X4 FILLER_87_926 ();
 FILLCELL_X2 FILLER_87_930 ();
 FILLCELL_X2 FILLER_87_938 ();
 FILLCELL_X4 FILLER_87_968 ();
 FILLCELL_X8 FILLER_87_993 ();
 FILLCELL_X4 FILLER_87_1001 ();
 FILLCELL_X1 FILLER_87_1005 ();
 FILLCELL_X16 FILLER_87_1016 ();
 FILLCELL_X8 FILLER_87_1032 ();
 FILLCELL_X2 FILLER_87_1040 ();
 FILLCELL_X2 FILLER_87_1060 ();
 FILLCELL_X1 FILLER_87_1062 ();
 FILLCELL_X2 FILLER_87_1067 ();
 FILLCELL_X8 FILLER_87_1082 ();
 FILLCELL_X1 FILLER_87_1090 ();
 FILLCELL_X4 FILLER_87_1096 ();
 FILLCELL_X2 FILLER_87_1100 ();
 FILLCELL_X1 FILLER_87_1102 ();
 FILLCELL_X1 FILLER_87_1106 ();
 FILLCELL_X4 FILLER_87_1118 ();
 FILLCELL_X2 FILLER_87_1122 ();
 FILLCELL_X1 FILLER_87_1124 ();
 FILLCELL_X2 FILLER_87_1132 ();
 FILLCELL_X8 FILLER_87_1141 ();
 FILLCELL_X4 FILLER_87_1149 ();
 FILLCELL_X2 FILLER_87_1153 ();
 FILLCELL_X1 FILLER_87_1159 ();
 FILLCELL_X1 FILLER_87_1172 ();
 FILLCELL_X1 FILLER_87_1177 ();
 FILLCELL_X8 FILLER_87_1189 ();
 FILLCELL_X2 FILLER_87_1197 ();
 FILLCELL_X1 FILLER_87_1199 ();
 FILLCELL_X4 FILLER_87_1203 ();
 FILLCELL_X2 FILLER_87_1207 ();
 FILLCELL_X16 FILLER_88_1 ();
 FILLCELL_X8 FILLER_88_17 ();
 FILLCELL_X2 FILLER_88_25 ();
 FILLCELL_X1 FILLER_88_27 ();
 FILLCELL_X32 FILLER_88_31 ();
 FILLCELL_X16 FILLER_88_63 ();
 FILLCELL_X4 FILLER_88_79 ();
 FILLCELL_X4 FILLER_88_94 ();
 FILLCELL_X2 FILLER_88_106 ();
 FILLCELL_X1 FILLER_88_108 ();
 FILLCELL_X2 FILLER_88_137 ();
 FILLCELL_X1 FILLER_88_139 ();
 FILLCELL_X2 FILLER_88_146 ();
 FILLCELL_X2 FILLER_88_162 ();
 FILLCELL_X1 FILLER_88_164 ();
 FILLCELL_X4 FILLER_88_188 ();
 FILLCELL_X16 FILLER_88_206 ();
 FILLCELL_X4 FILLER_88_222 ();
 FILLCELL_X2 FILLER_88_226 ();
 FILLCELL_X1 FILLER_88_228 ();
 FILLCELL_X4 FILLER_88_240 ();
 FILLCELL_X2 FILLER_88_244 ();
 FILLCELL_X1 FILLER_88_246 ();
 FILLCELL_X16 FILLER_88_256 ();
 FILLCELL_X4 FILLER_88_272 ();
 FILLCELL_X4 FILLER_88_293 ();
 FILLCELL_X2 FILLER_88_304 ();
 FILLCELL_X4 FILLER_88_316 ();
 FILLCELL_X2 FILLER_88_320 ();
 FILLCELL_X2 FILLER_88_339 ();
 FILLCELL_X2 FILLER_88_346 ();
 FILLCELL_X1 FILLER_88_348 ();
 FILLCELL_X1 FILLER_88_368 ();
 FILLCELL_X1 FILLER_88_375 ();
 FILLCELL_X2 FILLER_88_396 ();
 FILLCELL_X4 FILLER_88_407 ();
 FILLCELL_X1 FILLER_88_411 ();
 FILLCELL_X4 FILLER_88_436 ();
 FILLCELL_X2 FILLER_88_440 ();
 FILLCELL_X2 FILLER_88_448 ();
 FILLCELL_X16 FILLER_88_510 ();
 FILLCELL_X1 FILLER_88_526 ();
 FILLCELL_X2 FILLER_88_537 ();
 FILLCELL_X8 FILLER_88_544 ();
 FILLCELL_X2 FILLER_88_552 ();
 FILLCELL_X4 FILLER_88_569 ();
 FILLCELL_X16 FILLER_88_613 ();
 FILLCELL_X2 FILLER_88_629 ();
 FILLCELL_X8 FILLER_88_632 ();
 FILLCELL_X4 FILLER_88_640 ();
 FILLCELL_X2 FILLER_88_651 ();
 FILLCELL_X4 FILLER_88_671 ();
 FILLCELL_X2 FILLER_88_675 ();
 FILLCELL_X1 FILLER_88_681 ();
 FILLCELL_X1 FILLER_88_699 ();
 FILLCELL_X2 FILLER_88_719 ();
 FILLCELL_X1 FILLER_88_721 ();
 FILLCELL_X4 FILLER_88_739 ();
 FILLCELL_X16 FILLER_88_746 ();
 FILLCELL_X2 FILLER_88_762 ();
 FILLCELL_X1 FILLER_88_764 ();
 FILLCELL_X1 FILLER_88_802 ();
 FILLCELL_X1 FILLER_88_832 ();
 FILLCELL_X8 FILLER_88_839 ();
 FILLCELL_X4 FILLER_88_847 ();
 FILLCELL_X2 FILLER_88_851 ();
 FILLCELL_X4 FILLER_88_876 ();
 FILLCELL_X1 FILLER_88_889 ();
 FILLCELL_X2 FILLER_88_893 ();
 FILLCELL_X1 FILLER_88_895 ();
 FILLCELL_X8 FILLER_88_920 ();
 FILLCELL_X8 FILLER_88_940 ();
 FILLCELL_X2 FILLER_88_948 ();
 FILLCELL_X1 FILLER_88_950 ();
 FILLCELL_X1 FILLER_88_968 ();
 FILLCELL_X4 FILLER_88_1010 ();
 FILLCELL_X1 FILLER_88_1014 ();
 FILLCELL_X2 FILLER_88_1050 ();
 FILLCELL_X1 FILLER_88_1052 ();
 FILLCELL_X8 FILLER_88_1061 ();
 FILLCELL_X4 FILLER_88_1069 ();
 FILLCELL_X2 FILLER_88_1073 ();
 FILLCELL_X1 FILLER_88_1075 ();
 FILLCELL_X4 FILLER_88_1100 ();
 FILLCELL_X2 FILLER_88_1104 ();
 FILLCELL_X1 FILLER_88_1106 ();
 FILLCELL_X2 FILLER_88_1124 ();
 FILLCELL_X1 FILLER_88_1144 ();
 FILLCELL_X1 FILLER_88_1152 ();
 FILLCELL_X2 FILLER_88_1165 ();
 FILLCELL_X1 FILLER_88_1167 ();
 FILLCELL_X4 FILLER_88_1203 ();
 FILLCELL_X2 FILLER_88_1207 ();
 FILLCELL_X8 FILLER_89_4 ();
 FILLCELL_X2 FILLER_89_12 ();
 FILLCELL_X8 FILLER_89_21 ();
 FILLCELL_X1 FILLER_89_29 ();
 FILLCELL_X32 FILLER_89_33 ();
 FILLCELL_X16 FILLER_89_65 ();
 FILLCELL_X8 FILLER_89_81 ();
 FILLCELL_X2 FILLER_89_100 ();
 FILLCELL_X2 FILLER_89_108 ();
 FILLCELL_X2 FILLER_89_125 ();
 FILLCELL_X1 FILLER_89_127 ();
 FILLCELL_X1 FILLER_89_137 ();
 FILLCELL_X1 FILLER_89_142 ();
 FILLCELL_X8 FILLER_89_154 ();
 FILLCELL_X8 FILLER_89_168 ();
 FILLCELL_X2 FILLER_89_176 ();
 FILLCELL_X16 FILLER_89_191 ();
 FILLCELL_X8 FILLER_89_207 ();
 FILLCELL_X2 FILLER_89_215 ();
 FILLCELL_X8 FILLER_89_221 ();
 FILLCELL_X2 FILLER_89_229 ();
 FILLCELL_X1 FILLER_89_235 ();
 FILLCELL_X16 FILLER_89_241 ();
 FILLCELL_X4 FILLER_89_257 ();
 FILLCELL_X2 FILLER_89_261 ();
 FILLCELL_X4 FILLER_89_287 ();
 FILLCELL_X2 FILLER_89_296 ();
 FILLCELL_X2 FILLER_89_304 ();
 FILLCELL_X1 FILLER_89_306 ();
 FILLCELL_X8 FILLER_89_313 ();
 FILLCELL_X1 FILLER_89_321 ();
 FILLCELL_X1 FILLER_89_338 ();
 FILLCELL_X2 FILLER_89_345 ();
 FILLCELL_X1 FILLER_89_347 ();
 FILLCELL_X1 FILLER_89_352 ();
 FILLCELL_X8 FILLER_89_363 ();
 FILLCELL_X1 FILLER_89_371 ();
 FILLCELL_X8 FILLER_89_382 ();
 FILLCELL_X2 FILLER_89_390 ();
 FILLCELL_X8 FILLER_89_401 ();
 FILLCELL_X4 FILLER_89_409 ();
 FILLCELL_X2 FILLER_89_413 ();
 FILLCELL_X4 FILLER_89_436 ();
 FILLCELL_X4 FILLER_89_447 ();
 FILLCELL_X16 FILLER_89_460 ();
 FILLCELL_X1 FILLER_89_476 ();
 FILLCELL_X4 FILLER_89_507 ();
 FILLCELL_X2 FILLER_89_511 ();
 FILLCELL_X4 FILLER_89_520 ();
 FILLCELL_X2 FILLER_89_524 ();
 FILLCELL_X4 FILLER_89_533 ();
 FILLCELL_X1 FILLER_89_537 ();
 FILLCELL_X8 FILLER_89_542 ();
 FILLCELL_X2 FILLER_89_550 ();
 FILLCELL_X1 FILLER_89_556 ();
 FILLCELL_X16 FILLER_89_563 ();
 FILLCELL_X8 FILLER_89_579 ();
 FILLCELL_X1 FILLER_89_594 ();
 FILLCELL_X2 FILLER_89_598 ();
 FILLCELL_X8 FILLER_89_624 ();
 FILLCELL_X8 FILLER_89_639 ();
 FILLCELL_X2 FILLER_89_647 ();
 FILLCELL_X1 FILLER_89_649 ();
 FILLCELL_X32 FILLER_89_659 ();
 FILLCELL_X2 FILLER_89_691 ();
 FILLCELL_X1 FILLER_89_693 ();
 FILLCELL_X2 FILLER_89_711 ();
 FILLCELL_X1 FILLER_89_734 ();
 FILLCELL_X4 FILLER_89_738 ();
 FILLCELL_X1 FILLER_89_746 ();
 FILLCELL_X1 FILLER_89_753 ();
 FILLCELL_X8 FILLER_89_756 ();
 FILLCELL_X4 FILLER_89_764 ();
 FILLCELL_X2 FILLER_89_768 ();
 FILLCELL_X1 FILLER_89_770 ();
 FILLCELL_X4 FILLER_89_790 ();
 FILLCELL_X1 FILLER_89_794 ();
 FILLCELL_X1 FILLER_89_824 ();
 FILLCELL_X2 FILLER_89_853 ();
 FILLCELL_X1 FILLER_89_855 ();
 FILLCELL_X1 FILLER_89_866 ();
 FILLCELL_X8 FILLER_89_873 ();
 FILLCELL_X4 FILLER_89_881 ();
 FILLCELL_X1 FILLER_89_885 ();
 FILLCELL_X2 FILLER_89_899 ();
 FILLCELL_X2 FILLER_89_918 ();
 FILLCELL_X2 FILLER_89_930 ();
 FILLCELL_X1 FILLER_89_947 ();
 FILLCELL_X32 FILLER_89_954 ();
 FILLCELL_X2 FILLER_89_986 ();
 FILLCELL_X8 FILLER_89_1012 ();
 FILLCELL_X1 FILLER_89_1020 ();
 FILLCELL_X4 FILLER_89_1038 ();
 FILLCELL_X2 FILLER_89_1042 ();
 FILLCELL_X1 FILLER_89_1044 ();
 FILLCELL_X2 FILLER_89_1050 ();
 FILLCELL_X1 FILLER_89_1052 ();
 FILLCELL_X1 FILLER_89_1075 ();
 FILLCELL_X16 FILLER_89_1080 ();
 FILLCELL_X4 FILLER_89_1099 ();
 FILLCELL_X1 FILLER_89_1103 ();
 FILLCELL_X2 FILLER_89_1111 ();
 FILLCELL_X16 FILLER_89_1118 ();
 FILLCELL_X4 FILLER_89_1134 ();
 FILLCELL_X2 FILLER_89_1138 ();
 FILLCELL_X2 FILLER_89_1149 ();
 FILLCELL_X1 FILLER_89_1155 ();
 FILLCELL_X4 FILLER_89_1168 ();
 FILLCELL_X2 FILLER_89_1172 ();
 FILLCELL_X8 FILLER_89_1178 ();
 FILLCELL_X4 FILLER_89_1186 ();
 FILLCELL_X2 FILLER_89_1190 ();
 FILLCELL_X4 FILLER_89_1198 ();
 FILLCELL_X1 FILLER_89_1205 ();
 FILLCELL_X4 FILLER_90_1 ();
 FILLCELL_X2 FILLER_90_5 ();
 FILLCELL_X8 FILLER_90_10 ();
 FILLCELL_X4 FILLER_90_18 ();
 FILLCELL_X2 FILLER_90_22 ();
 FILLCELL_X1 FILLER_90_30 ();
 FILLCELL_X32 FILLER_90_34 ();
 FILLCELL_X16 FILLER_90_66 ();
 FILLCELL_X4 FILLER_90_82 ();
 FILLCELL_X4 FILLER_90_89 ();
 FILLCELL_X1 FILLER_90_97 ();
 FILLCELL_X2 FILLER_90_103 ();
 FILLCELL_X1 FILLER_90_105 ();
 FILLCELL_X4 FILLER_90_124 ();
 FILLCELL_X2 FILLER_90_128 ();
 FILLCELL_X2 FILLER_90_134 ();
 FILLCELL_X2 FILLER_90_140 ();
 FILLCELL_X8 FILLER_90_161 ();
 FILLCELL_X1 FILLER_90_174 ();
 FILLCELL_X4 FILLER_90_184 ();
 FILLCELL_X1 FILLER_90_188 ();
 FILLCELL_X4 FILLER_90_198 ();
 FILLCELL_X1 FILLER_90_202 ();
 FILLCELL_X2 FILLER_90_215 ();
 FILLCELL_X4 FILLER_90_220 ();
 FILLCELL_X2 FILLER_90_224 ();
 FILLCELL_X1 FILLER_90_226 ();
 FILLCELL_X2 FILLER_90_231 ();
 FILLCELL_X8 FILLER_90_240 ();
 FILLCELL_X1 FILLER_90_248 ();
 FILLCELL_X1 FILLER_90_266 ();
 FILLCELL_X4 FILLER_90_281 ();
 FILLCELL_X1 FILLER_90_285 ();
 FILLCELL_X2 FILLER_90_302 ();
 FILLCELL_X1 FILLER_90_304 ();
 FILLCELL_X4 FILLER_90_322 ();
 FILLCELL_X1 FILLER_90_396 ();
 FILLCELL_X8 FILLER_90_416 ();
 FILLCELL_X2 FILLER_90_439 ();
 FILLCELL_X32 FILLER_90_458 ();
 FILLCELL_X16 FILLER_90_490 ();
 FILLCELL_X4 FILLER_90_506 ();
 FILLCELL_X1 FILLER_90_510 ();
 FILLCELL_X1 FILLER_90_518 ();
 FILLCELL_X2 FILLER_90_529 ();
 FILLCELL_X2 FILLER_90_535 ();
 FILLCELL_X2 FILLER_90_544 ();
 FILLCELL_X4 FILLER_90_550 ();
 FILLCELL_X2 FILLER_90_554 ();
 FILLCELL_X1 FILLER_90_556 ();
 FILLCELL_X8 FILLER_90_568 ();
 FILLCELL_X1 FILLER_90_576 ();
 FILLCELL_X2 FILLER_90_584 ();
 FILLCELL_X1 FILLER_90_586 ();
 FILLCELL_X2 FILLER_90_591 ();
 FILLCELL_X1 FILLER_90_596 ();
 FILLCELL_X2 FILLER_90_612 ();
 FILLCELL_X8 FILLER_90_618 ();
 FILLCELL_X4 FILLER_90_626 ();
 FILLCELL_X1 FILLER_90_630 ();
 FILLCELL_X2 FILLER_90_632 ();
 FILLCELL_X1 FILLER_90_634 ();
 FILLCELL_X2 FILLER_90_655 ();
 FILLCELL_X1 FILLER_90_657 ();
 FILLCELL_X8 FILLER_90_665 ();
 FILLCELL_X1 FILLER_90_673 ();
 FILLCELL_X8 FILLER_90_752 ();
 FILLCELL_X4 FILLER_90_760 ();
 FILLCELL_X8 FILLER_90_780 ();
 FILLCELL_X2 FILLER_90_788 ();
 FILLCELL_X1 FILLER_90_790 ();
 FILLCELL_X1 FILLER_90_823 ();
 FILLCELL_X1 FILLER_90_837 ();
 FILLCELL_X8 FILLER_90_859 ();
 FILLCELL_X2 FILLER_90_887 ();
 FILLCELL_X8 FILLER_90_922 ();
 FILLCELL_X2 FILLER_90_936 ();
 FILLCELL_X1 FILLER_90_938 ();
 FILLCELL_X2 FILLER_90_945 ();
 FILLCELL_X1 FILLER_90_947 ();
 FILLCELL_X2 FILLER_90_989 ();
 FILLCELL_X1 FILLER_90_991 ();
 FILLCELL_X32 FILLER_90_996 ();
 FILLCELL_X16 FILLER_90_1028 ();
 FILLCELL_X4 FILLER_90_1044 ();
 FILLCELL_X2 FILLER_90_1048 ();
 FILLCELL_X1 FILLER_90_1050 ();
 FILLCELL_X2 FILLER_90_1083 ();
 FILLCELL_X2 FILLER_90_1088 ();
 FILLCELL_X4 FILLER_90_1108 ();
 FILLCELL_X2 FILLER_90_1112 ();
 FILLCELL_X1 FILLER_90_1129 ();
 FILLCELL_X2 FILLER_90_1153 ();
 FILLCELL_X2 FILLER_90_1167 ();
 FILLCELL_X8 FILLER_90_1180 ();
 FILLCELL_X2 FILLER_90_1188 ();
 FILLCELL_X1 FILLER_90_1190 ();
 FILLCELL_X8 FILLER_90_1194 ();
 FILLCELL_X4 FILLER_90_1202 ();
 FILLCELL_X2 FILLER_90_1206 ();
 FILLCELL_X1 FILLER_90_1208 ();
 FILLCELL_X2 FILLER_91_1 ();
 FILLCELL_X16 FILLER_91_9 ();
 FILLCELL_X4 FILLER_91_28 ();
 FILLCELL_X1 FILLER_91_32 ();
 FILLCELL_X32 FILLER_91_36 ();
 FILLCELL_X16 FILLER_91_68 ();
 FILLCELL_X4 FILLER_91_84 ();
 FILLCELL_X1 FILLER_91_104 ();
 FILLCELL_X2 FILLER_91_115 ();
 FILLCELL_X2 FILLER_91_125 ();
 FILLCELL_X1 FILLER_91_127 ();
 FILLCELL_X1 FILLER_91_132 ();
 FILLCELL_X1 FILLER_91_137 ();
 FILLCELL_X8 FILLER_91_151 ();
 FILLCELL_X4 FILLER_91_159 ();
 FILLCELL_X2 FILLER_91_163 ();
 FILLCELL_X1 FILLER_91_165 ();
 FILLCELL_X1 FILLER_91_183 ();
 FILLCELL_X2 FILLER_91_188 ();
 FILLCELL_X1 FILLER_91_206 ();
 FILLCELL_X2 FILLER_91_222 ();
 FILLCELL_X2 FILLER_91_240 ();
 FILLCELL_X1 FILLER_91_242 ();
 FILLCELL_X1 FILLER_91_250 ();
 FILLCELL_X2 FILLER_91_268 ();
 FILLCELL_X1 FILLER_91_287 ();
 FILLCELL_X2 FILLER_91_303 ();
 FILLCELL_X4 FILLER_91_312 ();
 FILLCELL_X1 FILLER_91_316 ();
 FILLCELL_X2 FILLER_91_339 ();
 FILLCELL_X4 FILLER_91_348 ();
 FILLCELL_X1 FILLER_91_352 ();
 FILLCELL_X4 FILLER_91_356 ();
 FILLCELL_X1 FILLER_91_363 ();
 FILLCELL_X2 FILLER_91_390 ();
 FILLCELL_X4 FILLER_91_420 ();
 FILLCELL_X2 FILLER_91_424 ();
 FILLCELL_X8 FILLER_91_443 ();
 FILLCELL_X2 FILLER_91_451 ();
 FILLCELL_X4 FILLER_91_466 ();
 FILLCELL_X2 FILLER_91_470 ();
 FILLCELL_X8 FILLER_91_489 ();
 FILLCELL_X4 FILLER_91_497 ();
 FILLCELL_X2 FILLER_91_501 ();
 FILLCELL_X1 FILLER_91_503 ();
 FILLCELL_X8 FILLER_91_509 ();
 FILLCELL_X4 FILLER_91_517 ();
 FILLCELL_X1 FILLER_91_521 ();
 FILLCELL_X4 FILLER_91_528 ();
 FILLCELL_X1 FILLER_91_532 ();
 FILLCELL_X4 FILLER_91_536 ();
 FILLCELL_X2 FILLER_91_546 ();
 FILLCELL_X1 FILLER_91_548 ();
 FILLCELL_X32 FILLER_91_553 ();
 FILLCELL_X16 FILLER_91_603 ();
 FILLCELL_X8 FILLER_91_619 ();
 FILLCELL_X2 FILLER_91_635 ();
 FILLCELL_X2 FILLER_91_641 ();
 FILLCELL_X2 FILLER_91_662 ();
 FILLCELL_X1 FILLER_91_664 ();
 FILLCELL_X16 FILLER_91_669 ();
 FILLCELL_X8 FILLER_91_685 ();
 FILLCELL_X4 FILLER_91_693 ();
 FILLCELL_X2 FILLER_91_697 ();
 FILLCELL_X8 FILLER_91_704 ();
 FILLCELL_X4 FILLER_91_712 ();
 FILLCELL_X2 FILLER_91_716 ();
 FILLCELL_X2 FILLER_91_739 ();
 FILLCELL_X2 FILLER_91_769 ();
 FILLCELL_X1 FILLER_91_771 ();
 FILLCELL_X1 FILLER_91_785 ();
 FILLCELL_X1 FILLER_91_791 ();
 FILLCELL_X1 FILLER_91_812 ();
 FILLCELL_X4 FILLER_91_832 ();
 FILLCELL_X2 FILLER_91_836 ();
 FILLCELL_X16 FILLER_91_848 ();
 FILLCELL_X4 FILLER_91_864 ();
 FILLCELL_X2 FILLER_91_887 ();
 FILLCELL_X2 FILLER_91_896 ();
 FILLCELL_X8 FILLER_91_928 ();
 FILLCELL_X1 FILLER_91_942 ();
 FILLCELL_X8 FILLER_91_949 ();
 FILLCELL_X4 FILLER_91_957 ();
 FILLCELL_X1 FILLER_91_961 ();
 FILLCELL_X2 FILLER_91_971 ();
 FILLCELL_X1 FILLER_91_997 ();
 FILLCELL_X8 FILLER_91_1005 ();
 FILLCELL_X16 FILLER_91_1019 ();
 FILLCELL_X4 FILLER_91_1035 ();
 FILLCELL_X2 FILLER_91_1039 ();
 FILLCELL_X32 FILLER_91_1058 ();
 FILLCELL_X4 FILLER_91_1090 ();
 FILLCELL_X2 FILLER_91_1094 ();
 FILLCELL_X32 FILLER_91_1100 ();
 FILLCELL_X32 FILLER_91_1132 ();
 FILLCELL_X8 FILLER_91_1164 ();
 FILLCELL_X2 FILLER_91_1172 ();
 FILLCELL_X1 FILLER_91_1174 ();
 FILLCELL_X4 FILLER_91_1178 ();
 FILLCELL_X2 FILLER_91_1182 ();
 FILLCELL_X8 FILLER_91_1187 ();
 FILLCELL_X1 FILLER_91_1195 ();
 FILLCELL_X1 FILLER_91_1199 ();
 FILLCELL_X2 FILLER_91_1203 ();
 FILLCELL_X4 FILLER_92_1 ();
 FILLCELL_X2 FILLER_92_5 ();
 FILLCELL_X16 FILLER_92_10 ();
 FILLCELL_X2 FILLER_92_26 ();
 FILLCELL_X32 FILLER_92_31 ();
 FILLCELL_X32 FILLER_92_63 ();
 FILLCELL_X8 FILLER_92_95 ();
 FILLCELL_X4 FILLER_92_103 ();
 FILLCELL_X2 FILLER_92_107 ();
 FILLCELL_X1 FILLER_92_109 ();
 FILLCELL_X2 FILLER_92_114 ();
 FILLCELL_X8 FILLER_92_125 ();
 FILLCELL_X4 FILLER_92_133 ();
 FILLCELL_X2 FILLER_92_137 ();
 FILLCELL_X1 FILLER_92_139 ();
 FILLCELL_X2 FILLER_92_146 ();
 FILLCELL_X1 FILLER_92_148 ();
 FILLCELL_X1 FILLER_92_152 ();
 FILLCELL_X2 FILLER_92_157 ();
 FILLCELL_X2 FILLER_92_163 ();
 FILLCELL_X8 FILLER_92_170 ();
 FILLCELL_X1 FILLER_92_195 ();
 FILLCELL_X4 FILLER_92_204 ();
 FILLCELL_X2 FILLER_92_212 ();
 FILLCELL_X1 FILLER_92_214 ();
 FILLCELL_X32 FILLER_92_238 ();
 FILLCELL_X2 FILLER_92_270 ();
 FILLCELL_X1 FILLER_92_272 ();
 FILLCELL_X1 FILLER_92_289 ();
 FILLCELL_X8 FILLER_92_304 ();
 FILLCELL_X4 FILLER_92_312 ();
 FILLCELL_X2 FILLER_92_316 ();
 FILLCELL_X4 FILLER_92_339 ();
 FILLCELL_X1 FILLER_92_343 ();
 FILLCELL_X2 FILLER_92_363 ();
 FILLCELL_X1 FILLER_92_385 ();
 FILLCELL_X4 FILLER_92_390 ();
 FILLCELL_X4 FILLER_92_422 ();
 FILLCELL_X1 FILLER_92_426 ();
 FILLCELL_X8 FILLER_92_436 ();
 FILLCELL_X1 FILLER_92_444 ();
 FILLCELL_X4 FILLER_92_452 ();
 FILLCELL_X2 FILLER_92_456 ();
 FILLCELL_X1 FILLER_92_458 ();
 FILLCELL_X16 FILLER_92_493 ();
 FILLCELL_X4 FILLER_92_509 ();
 FILLCELL_X1 FILLER_92_513 ();
 FILLCELL_X4 FILLER_92_521 ();
 FILLCELL_X2 FILLER_92_525 ();
 FILLCELL_X2 FILLER_92_558 ();
 FILLCELL_X2 FILLER_92_563 ();
 FILLCELL_X1 FILLER_92_575 ();
 FILLCELL_X2 FILLER_92_583 ();
 FILLCELL_X1 FILLER_92_585 ();
 FILLCELL_X4 FILLER_92_611 ();
 FILLCELL_X2 FILLER_92_615 ();
 FILLCELL_X2 FILLER_92_628 ();
 FILLCELL_X1 FILLER_92_630 ();
 FILLCELL_X2 FILLER_92_646 ();
 FILLCELL_X1 FILLER_92_648 ();
 FILLCELL_X16 FILLER_92_667 ();
 FILLCELL_X2 FILLER_92_683 ();
 FILLCELL_X4 FILLER_92_711 ();
 FILLCELL_X2 FILLER_92_715 ();
 FILLCELL_X1 FILLER_92_717 ();
 FILLCELL_X2 FILLER_92_721 ();
 FILLCELL_X1 FILLER_92_723 ();
 FILLCELL_X16 FILLER_92_733 ();
 FILLCELL_X1 FILLER_92_749 ();
 FILLCELL_X4 FILLER_92_771 ();
 FILLCELL_X1 FILLER_92_775 ();
 FILLCELL_X4 FILLER_92_797 ();
 FILLCELL_X2 FILLER_92_813 ();
 FILLCELL_X2 FILLER_92_830 ();
 FILLCELL_X1 FILLER_92_892 ();
 FILLCELL_X8 FILLER_92_911 ();
 FILLCELL_X4 FILLER_92_940 ();
 FILLCELL_X2 FILLER_92_944 ();
 FILLCELL_X1 FILLER_92_946 ();
 FILLCELL_X2 FILLER_92_962 ();
 FILLCELL_X8 FILLER_92_967 ();
 FILLCELL_X1 FILLER_92_975 ();
 FILLCELL_X8 FILLER_92_1009 ();
 FILLCELL_X32 FILLER_92_1036 ();
 FILLCELL_X16 FILLER_92_1068 ();
 FILLCELL_X8 FILLER_92_1084 ();
 FILLCELL_X32 FILLER_92_1103 ();
 FILLCELL_X32 FILLER_92_1135 ();
 FILLCELL_X32 FILLER_92_1167 ();
 FILLCELL_X2 FILLER_92_1199 ();
 FILLCELL_X1 FILLER_92_1204 ();
 FILLCELL_X8 FILLER_93_1 ();
 FILLCELL_X4 FILLER_93_9 ();
 FILLCELL_X32 FILLER_93_16 ();
 FILLCELL_X32 FILLER_93_48 ();
 FILLCELL_X16 FILLER_93_80 ();
 FILLCELL_X8 FILLER_93_96 ();
 FILLCELL_X1 FILLER_93_104 ();
 FILLCELL_X8 FILLER_93_115 ();
 FILLCELL_X1 FILLER_93_123 ();
 FILLCELL_X1 FILLER_93_136 ();
 FILLCELL_X4 FILLER_93_144 ();
 FILLCELL_X2 FILLER_93_148 ();
 FILLCELL_X4 FILLER_93_154 ();
 FILLCELL_X2 FILLER_93_158 ();
 FILLCELL_X1 FILLER_93_166 ();
 FILLCELL_X16 FILLER_93_177 ();
 FILLCELL_X8 FILLER_93_193 ();
 FILLCELL_X4 FILLER_93_201 ();
 FILLCELL_X2 FILLER_93_205 ();
 FILLCELL_X1 FILLER_93_207 ();
 FILLCELL_X8 FILLER_93_215 ();
 FILLCELL_X4 FILLER_93_223 ();
 FILLCELL_X1 FILLER_93_227 ();
 FILLCELL_X16 FILLER_93_232 ();
 FILLCELL_X1 FILLER_93_265 ();
 FILLCELL_X2 FILLER_93_285 ();
 FILLCELL_X1 FILLER_93_295 ();
 FILLCELL_X16 FILLER_93_306 ();
 FILLCELL_X4 FILLER_93_322 ();
 FILLCELL_X4 FILLER_93_352 ();
 FILLCELL_X2 FILLER_93_356 ();
 FILLCELL_X1 FILLER_93_358 ();
 FILLCELL_X8 FILLER_93_362 ();
 FILLCELL_X4 FILLER_93_370 ();
 FILLCELL_X1 FILLER_93_374 ();
 FILLCELL_X4 FILLER_93_388 ();
 FILLCELL_X1 FILLER_93_396 ();
 FILLCELL_X1 FILLER_93_400 ();
 FILLCELL_X1 FILLER_93_408 ();
 FILLCELL_X2 FILLER_93_412 ();
 FILLCELL_X32 FILLER_93_417 ();
 FILLCELL_X4 FILLER_93_449 ();
 FILLCELL_X2 FILLER_93_453 ();
 FILLCELL_X8 FILLER_93_462 ();
 FILLCELL_X4 FILLER_93_470 ();
 FILLCELL_X1 FILLER_93_474 ();
 FILLCELL_X16 FILLER_93_489 ();
 FILLCELL_X8 FILLER_93_505 ();
 FILLCELL_X2 FILLER_93_513 ();
 FILLCELL_X2 FILLER_93_519 ();
 FILLCELL_X1 FILLER_93_521 ();
 FILLCELL_X4 FILLER_93_532 ();
 FILLCELL_X8 FILLER_93_542 ();
 FILLCELL_X1 FILLER_93_550 ();
 FILLCELL_X2 FILLER_93_560 ();
 FILLCELL_X8 FILLER_93_566 ();
 FILLCELL_X1 FILLER_93_574 ();
 FILLCELL_X1 FILLER_93_582 ();
 FILLCELL_X4 FILLER_93_606 ();
 FILLCELL_X1 FILLER_93_610 ();
 FILLCELL_X4 FILLER_93_617 ();
 FILLCELL_X2 FILLER_93_621 ();
 FILLCELL_X4 FILLER_93_649 ();
 FILLCELL_X32 FILLER_93_659 ();
 FILLCELL_X16 FILLER_93_691 ();
 FILLCELL_X8 FILLER_93_707 ();
 FILLCELL_X4 FILLER_93_715 ();
 FILLCELL_X4 FILLER_93_735 ();
 FILLCELL_X2 FILLER_93_739 ();
 FILLCELL_X8 FILLER_93_748 ();
 FILLCELL_X4 FILLER_93_756 ();
 FILLCELL_X1 FILLER_93_760 ();
 FILLCELL_X2 FILLER_93_782 ();
 FILLCELL_X1 FILLER_93_795 ();
 FILLCELL_X8 FILLER_93_811 ();
 FILLCELL_X2 FILLER_93_819 ();
 FILLCELL_X1 FILLER_93_840 ();
 FILLCELL_X1 FILLER_93_844 ();
 FILLCELL_X8 FILLER_93_855 ();
 FILLCELL_X4 FILLER_93_863 ();
 FILLCELL_X1 FILLER_93_873 ();
 FILLCELL_X1 FILLER_93_906 ();
 FILLCELL_X8 FILLER_93_940 ();
 FILLCELL_X2 FILLER_93_948 ();
 FILLCELL_X2 FILLER_93_953 ();
 FILLCELL_X1 FILLER_93_955 ();
 FILLCELL_X1 FILLER_93_958 ();
 FILLCELL_X1 FILLER_93_962 ();
 FILLCELL_X8 FILLER_93_972 ();
 FILLCELL_X2 FILLER_93_994 ();
 FILLCELL_X1 FILLER_93_996 ();
 FILLCELL_X16 FILLER_93_1003 ();
 FILLCELL_X8 FILLER_93_1019 ();
 FILLCELL_X4 FILLER_93_1034 ();
 FILLCELL_X2 FILLER_93_1038 ();
 FILLCELL_X1 FILLER_93_1040 ();
 FILLCELL_X16 FILLER_93_1058 ();
 FILLCELL_X8 FILLER_93_1074 ();
 FILLCELL_X2 FILLER_93_1082 ();
 FILLCELL_X32 FILLER_93_1101 ();
 FILLCELL_X32 FILLER_93_1133 ();
 FILLCELL_X4 FILLER_93_1165 ();
 FILLCELL_X1 FILLER_93_1169 ();
 FILLCELL_X8 FILLER_93_1173 ();
 FILLCELL_X2 FILLER_93_1181 ();
 FILLCELL_X1 FILLER_93_1183 ();
 FILLCELL_X4 FILLER_93_1187 ();
 FILLCELL_X8 FILLER_93_1194 ();
 FILLCELL_X2 FILLER_93_1202 ();
 FILLCELL_X1 FILLER_93_1204 ();
 FILLCELL_X16 FILLER_94_4 ();
 FILLCELL_X2 FILLER_94_20 ();
 FILLCELL_X2 FILLER_94_25 ();
 FILLCELL_X4 FILLER_94_31 ();
 FILLCELL_X2 FILLER_94_35 ();
 FILLCELL_X32 FILLER_94_40 ();
 FILLCELL_X32 FILLER_94_72 ();
 FILLCELL_X32 FILLER_94_104 ();
 FILLCELL_X16 FILLER_94_136 ();
 FILLCELL_X4 FILLER_94_152 ();
 FILLCELL_X8 FILLER_94_163 ();
 FILLCELL_X4 FILLER_94_171 ();
 FILLCELL_X16 FILLER_94_182 ();
 FILLCELL_X8 FILLER_94_198 ();
 FILLCELL_X2 FILLER_94_206 ();
 FILLCELL_X1 FILLER_94_208 ();
 FILLCELL_X16 FILLER_94_250 ();
 FILLCELL_X8 FILLER_94_266 ();
 FILLCELL_X2 FILLER_94_284 ();
 FILLCELL_X4 FILLER_94_290 ();
 FILLCELL_X2 FILLER_94_294 ();
 FILLCELL_X2 FILLER_94_302 ();
 FILLCELL_X1 FILLER_94_304 ();
 FILLCELL_X2 FILLER_94_329 ();
 FILLCELL_X4 FILLER_94_347 ();
 FILLCELL_X2 FILLER_94_351 ();
 FILLCELL_X2 FILLER_94_387 ();
 FILLCELL_X1 FILLER_94_399 ();
 FILLCELL_X2 FILLER_94_404 ();
 FILLCELL_X1 FILLER_94_419 ();
 FILLCELL_X16 FILLER_94_427 ();
 FILLCELL_X2 FILLER_94_443 ();
 FILLCELL_X4 FILLER_94_452 ();
 FILLCELL_X4 FILLER_94_464 ();
 FILLCELL_X32 FILLER_94_475 ();
 FILLCELL_X2 FILLER_94_507 ();
 FILLCELL_X4 FILLER_94_519 ();
 FILLCELL_X1 FILLER_94_523 ();
 FILLCELL_X8 FILLER_94_529 ();
 FILLCELL_X2 FILLER_94_537 ();
 FILLCELL_X2 FILLER_94_550 ();
 FILLCELL_X4 FILLER_94_567 ();
 FILLCELL_X2 FILLER_94_571 ();
 FILLCELL_X1 FILLER_94_573 ();
 FILLCELL_X4 FILLER_94_587 ();
 FILLCELL_X1 FILLER_94_602 ();
 FILLCELL_X2 FILLER_94_608 ();
 FILLCELL_X1 FILLER_94_610 ();
 FILLCELL_X8 FILLER_94_618 ();
 FILLCELL_X1 FILLER_94_626 ();
 FILLCELL_X2 FILLER_94_632 ();
 FILLCELL_X1 FILLER_94_634 ();
 FILLCELL_X8 FILLER_94_638 ();
 FILLCELL_X2 FILLER_94_649 ();
 FILLCELL_X1 FILLER_94_651 ();
 FILLCELL_X32 FILLER_94_656 ();
 FILLCELL_X8 FILLER_94_714 ();
 FILLCELL_X1 FILLER_94_729 ();
 FILLCELL_X4 FILLER_94_743 ();
 FILLCELL_X2 FILLER_94_747 ();
 FILLCELL_X1 FILLER_94_749 ();
 FILLCELL_X1 FILLER_94_805 ();
 FILLCELL_X2 FILLER_94_815 ();
 FILLCELL_X1 FILLER_94_817 ();
 FILLCELL_X1 FILLER_94_834 ();
 FILLCELL_X8 FILLER_94_851 ();
 FILLCELL_X1 FILLER_94_859 ();
 FILLCELL_X2 FILLER_94_869 ();
 FILLCELL_X8 FILLER_94_907 ();
 FILLCELL_X4 FILLER_94_919 ();
 FILLCELL_X1 FILLER_94_923 ();
 FILLCELL_X4 FILLER_94_935 ();
 FILLCELL_X2 FILLER_94_939 ();
 FILLCELL_X1 FILLER_94_941 ();
 FILLCELL_X4 FILLER_94_972 ();
 FILLCELL_X2 FILLER_94_976 ();
 FILLCELL_X1 FILLER_94_978 ();
 FILLCELL_X4 FILLER_94_986 ();
 FILLCELL_X2 FILLER_94_990 ();
 FILLCELL_X1 FILLER_94_1001 ();
 FILLCELL_X1 FILLER_94_1019 ();
 FILLCELL_X16 FILLER_94_1029 ();
 FILLCELL_X8 FILLER_94_1045 ();
 FILLCELL_X16 FILLER_94_1062 ();
 FILLCELL_X4 FILLER_94_1078 ();
 FILLCELL_X2 FILLER_94_1082 ();
 FILLCELL_X1 FILLER_94_1084 ();
 FILLCELL_X1 FILLER_94_1102 ();
 FILLCELL_X8 FILLER_94_1122 ();
 FILLCELL_X2 FILLER_94_1130 ();
 FILLCELL_X32 FILLER_94_1156 ();
 FILLCELL_X1 FILLER_94_1191 ();
 FILLCELL_X8 FILLER_94_1195 ();
 FILLCELL_X4 FILLER_94_1203 ();
 FILLCELL_X2 FILLER_94_1207 ();
 FILLCELL_X2 FILLER_95_1 ();
 FILLCELL_X8 FILLER_95_6 ();
 FILLCELL_X8 FILLER_95_21 ();
 FILLCELL_X2 FILLER_95_29 ();
 FILLCELL_X1 FILLER_95_31 ();
 FILLCELL_X32 FILLER_95_35 ();
 FILLCELL_X32 FILLER_95_67 ();
 FILLCELL_X32 FILLER_95_99 ();
 FILLCELL_X16 FILLER_95_131 ();
 FILLCELL_X8 FILLER_95_147 ();
 FILLCELL_X1 FILLER_95_155 ();
 FILLCELL_X32 FILLER_95_192 ();
 FILLCELL_X8 FILLER_95_224 ();
 FILLCELL_X16 FILLER_95_239 ();
 FILLCELL_X2 FILLER_95_255 ();
 FILLCELL_X1 FILLER_95_257 ();
 FILLCELL_X2 FILLER_95_283 ();
 FILLCELL_X1 FILLER_95_285 ();
 FILLCELL_X8 FILLER_95_312 ();
 FILLCELL_X4 FILLER_95_320 ();
 FILLCELL_X2 FILLER_95_324 ();
 FILLCELL_X1 FILLER_95_326 ();
 FILLCELL_X4 FILLER_95_333 ();
 FILLCELL_X4 FILLER_95_384 ();
 FILLCELL_X1 FILLER_95_394 ();
 FILLCELL_X1 FILLER_95_406 ();
 FILLCELL_X2 FILLER_95_424 ();
 FILLCELL_X8 FILLER_95_437 ();
 FILLCELL_X4 FILLER_95_445 ();
 FILLCELL_X2 FILLER_95_449 ();
 FILLCELL_X1 FILLER_95_451 ();
 FILLCELL_X16 FILLER_95_482 ();
 FILLCELL_X8 FILLER_95_498 ();
 FILLCELL_X1 FILLER_95_506 ();
 FILLCELL_X4 FILLER_95_510 ();
 FILLCELL_X2 FILLER_95_514 ();
 FILLCELL_X1 FILLER_95_516 ();
 FILLCELL_X2 FILLER_95_520 ();
 FILLCELL_X8 FILLER_95_559 ();
 FILLCELL_X4 FILLER_95_567 ();
 FILLCELL_X2 FILLER_95_571 ();
 FILLCELL_X1 FILLER_95_573 ();
 FILLCELL_X16 FILLER_95_586 ();
 FILLCELL_X2 FILLER_95_602 ();
 FILLCELL_X1 FILLER_95_616 ();
 FILLCELL_X1 FILLER_95_624 ();
 FILLCELL_X4 FILLER_95_632 ();
 FILLCELL_X2 FILLER_95_636 ();
 FILLCELL_X4 FILLER_95_652 ();
 FILLCELL_X2 FILLER_95_656 ();
 FILLCELL_X4 FILLER_95_675 ();
 FILLCELL_X2 FILLER_95_679 ();
 FILLCELL_X1 FILLER_95_681 ();
 FILLCELL_X16 FILLER_95_703 ();
 FILLCELL_X4 FILLER_95_719 ();
 FILLCELL_X1 FILLER_95_729 ();
 FILLCELL_X8 FILLER_95_737 ();
 FILLCELL_X4 FILLER_95_745 ();
 FILLCELL_X2 FILLER_95_771 ();
 FILLCELL_X2 FILLER_95_802 ();
 FILLCELL_X4 FILLER_95_814 ();
 FILLCELL_X2 FILLER_95_818 ();
 FILLCELL_X1 FILLER_95_820 ();
 FILLCELL_X2 FILLER_95_824 ();
 FILLCELL_X1 FILLER_95_826 ();
 FILLCELL_X1 FILLER_95_901 ();
 FILLCELL_X16 FILLER_95_912 ();
 FILLCELL_X4 FILLER_95_928 ();
 FILLCELL_X2 FILLER_95_932 ();
 FILLCELL_X1 FILLER_95_934 ();
 FILLCELL_X8 FILLER_95_996 ();
 FILLCELL_X4 FILLER_95_1004 ();
 FILLCELL_X2 FILLER_95_1008 ();
 FILLCELL_X1 FILLER_95_1010 ();
 FILLCELL_X8 FILLER_95_1030 ();
 FILLCELL_X4 FILLER_95_1038 ();
 FILLCELL_X4 FILLER_95_1063 ();
 FILLCELL_X1 FILLER_95_1067 ();
 FILLCELL_X1 FILLER_95_1075 ();
 FILLCELL_X1 FILLER_95_1085 ();
 FILLCELL_X2 FILLER_95_1102 ();
 FILLCELL_X16 FILLER_95_1125 ();
 FILLCELL_X8 FILLER_95_1141 ();
 FILLCELL_X1 FILLER_95_1149 ();
 FILLCELL_X1 FILLER_95_1181 ();
 FILLCELL_X16 FILLER_95_1185 ();
 FILLCELL_X8 FILLER_95_1201 ();
 FILLCELL_X32 FILLER_96_1 ();
 FILLCELL_X2 FILLER_96_33 ();
 FILLCELL_X32 FILLER_96_38 ();
 FILLCELL_X32 FILLER_96_70 ();
 FILLCELL_X16 FILLER_96_102 ();
 FILLCELL_X8 FILLER_96_118 ();
 FILLCELL_X4 FILLER_96_126 ();
 FILLCELL_X2 FILLER_96_130 ();
 FILLCELL_X32 FILLER_96_149 ();
 FILLCELL_X32 FILLER_96_181 ();
 FILLCELL_X2 FILLER_96_213 ();
 FILLCELL_X1 FILLER_96_215 ();
 FILLCELL_X4 FILLER_96_238 ();
 FILLCELL_X2 FILLER_96_242 ();
 FILLCELL_X1 FILLER_96_244 ();
 FILLCELL_X2 FILLER_96_267 ();
 FILLCELL_X1 FILLER_96_284 ();
 FILLCELL_X4 FILLER_96_298 ();
 FILLCELL_X2 FILLER_96_306 ();
 FILLCELL_X1 FILLER_96_308 ();
 FILLCELL_X4 FILLER_96_318 ();
 FILLCELL_X2 FILLER_96_322 ();
 FILLCELL_X1 FILLER_96_324 ();
 FILLCELL_X4 FILLER_96_332 ();
 FILLCELL_X1 FILLER_96_336 ();
 FILLCELL_X1 FILLER_96_358 ();
 FILLCELL_X4 FILLER_96_362 ();
 FILLCELL_X2 FILLER_96_366 ();
 FILLCELL_X1 FILLER_96_368 ();
 FILLCELL_X2 FILLER_96_379 ();
 FILLCELL_X1 FILLER_96_381 ();
 FILLCELL_X4 FILLER_96_402 ();
 FILLCELL_X1 FILLER_96_406 ();
 FILLCELL_X32 FILLER_96_410 ();
 FILLCELL_X16 FILLER_96_442 ();
 FILLCELL_X16 FILLER_96_487 ();
 FILLCELL_X1 FILLER_96_503 ();
 FILLCELL_X4 FILLER_96_511 ();
 FILLCELL_X2 FILLER_96_515 ();
 FILLCELL_X8 FILLER_96_524 ();
 FILLCELL_X4 FILLER_96_532 ();
 FILLCELL_X2 FILLER_96_536 ();
 FILLCELL_X1 FILLER_96_538 ();
 FILLCELL_X2 FILLER_96_542 ();
 FILLCELL_X1 FILLER_96_544 ();
 FILLCELL_X8 FILLER_96_555 ();
 FILLCELL_X8 FILLER_96_570 ();
 FILLCELL_X1 FILLER_96_578 ();
 FILLCELL_X16 FILLER_96_586 ();
 FILLCELL_X16 FILLER_96_609 ();
 FILLCELL_X1 FILLER_96_625 ();
 FILLCELL_X4 FILLER_96_632 ();
 FILLCELL_X2 FILLER_96_636 ();
 FILLCELL_X1 FILLER_96_638 ();
 FILLCELL_X4 FILLER_96_643 ();
 FILLCELL_X2 FILLER_96_647 ();
 FILLCELL_X1 FILLER_96_649 ();
 FILLCELL_X2 FILLER_96_655 ();
 FILLCELL_X8 FILLER_96_661 ();
 FILLCELL_X2 FILLER_96_669 ();
 FILLCELL_X1 FILLER_96_671 ();
 FILLCELL_X1 FILLER_96_683 ();
 FILLCELL_X8 FILLER_96_707 ();
 FILLCELL_X2 FILLER_96_715 ();
 FILLCELL_X1 FILLER_96_717 ();
 FILLCELL_X4 FILLER_96_744 ();
 FILLCELL_X1 FILLER_96_748 ();
 FILLCELL_X2 FILLER_96_759 ();
 FILLCELL_X1 FILLER_96_764 ();
 FILLCELL_X1 FILLER_96_769 ();
 FILLCELL_X2 FILLER_96_784 ();
 FILLCELL_X2 FILLER_96_816 ();
 FILLCELL_X8 FILLER_96_825 ();
 FILLCELL_X1 FILLER_96_833 ();
 FILLCELL_X1 FILLER_96_848 ();
 FILLCELL_X2 FILLER_96_856 ();
 FILLCELL_X1 FILLER_96_871 ();
 FILLCELL_X2 FILLER_96_878 ();
 FILLCELL_X4 FILLER_96_883 ();
 FILLCELL_X2 FILLER_96_887 ();
 FILLCELL_X8 FILLER_96_892 ();
 FILLCELL_X2 FILLER_96_900 ();
 FILLCELL_X1 FILLER_96_902 ();
 FILLCELL_X4 FILLER_96_908 ();
 FILLCELL_X1 FILLER_96_912 ();
 FILLCELL_X4 FILLER_96_928 ();
 FILLCELL_X2 FILLER_96_932 ();
 FILLCELL_X2 FILLER_96_947 ();
 FILLCELL_X1 FILLER_96_971 ();
 FILLCELL_X8 FILLER_96_978 ();
 FILLCELL_X4 FILLER_96_986 ();
 FILLCELL_X2 FILLER_96_990 ();
 FILLCELL_X1 FILLER_96_992 ();
 FILLCELL_X16 FILLER_96_1010 ();
 FILLCELL_X2 FILLER_96_1026 ();
 FILLCELL_X4 FILLER_96_1035 ();
 FILLCELL_X2 FILLER_96_1039 ();
 FILLCELL_X1 FILLER_96_1041 ();
 FILLCELL_X8 FILLER_96_1074 ();
 FILLCELL_X4 FILLER_96_1082 ();
 FILLCELL_X4 FILLER_96_1106 ();
 FILLCELL_X2 FILLER_96_1110 ();
 FILLCELL_X1 FILLER_96_1136 ();
 FILLCELL_X4 FILLER_96_1142 ();
 FILLCELL_X1 FILLER_96_1146 ();
 FILLCELL_X2 FILLER_96_1162 ();
 FILLCELL_X1 FILLER_96_1164 ();
 FILLCELL_X2 FILLER_96_1182 ();
 FILLCELL_X1 FILLER_96_1184 ();
 FILLCELL_X1 FILLER_96_1188 ();
 FILLCELL_X4 FILLER_96_1198 ();
 FILLCELL_X2 FILLER_96_1206 ();
 FILLCELL_X1 FILLER_96_1208 ();
 FILLCELL_X4 FILLER_97_1 ();
 FILLCELL_X2 FILLER_97_5 ();
 FILLCELL_X32 FILLER_97_10 ();
 FILLCELL_X32 FILLER_97_42 ();
 FILLCELL_X32 FILLER_97_74 ();
 FILLCELL_X8 FILLER_97_106 ();
 FILLCELL_X2 FILLER_97_114 ();
 FILLCELL_X1 FILLER_97_116 ();
 FILLCELL_X4 FILLER_97_124 ();
 FILLCELL_X2 FILLER_97_128 ();
 FILLCELL_X1 FILLER_97_130 ();
 FILLCELL_X4 FILLER_97_151 ();
 FILLCELL_X2 FILLER_97_155 ();
 FILLCELL_X1 FILLER_97_157 ();
 FILLCELL_X2 FILLER_97_188 ();
 FILLCELL_X2 FILLER_97_226 ();
 FILLCELL_X2 FILLER_97_262 ();
 FILLCELL_X2 FILLER_97_284 ();
 FILLCELL_X4 FILLER_97_293 ();
 FILLCELL_X2 FILLER_97_297 ();
 FILLCELL_X1 FILLER_97_299 ();
 FILLCELL_X4 FILLER_97_320 ();
 FILLCELL_X2 FILLER_97_324 ();
 FILLCELL_X1 FILLER_97_326 ();
 FILLCELL_X4 FILLER_97_337 ();
 FILLCELL_X1 FILLER_97_359 ();
 FILLCELL_X4 FILLER_97_363 ();
 FILLCELL_X2 FILLER_97_367 ();
 FILLCELL_X1 FILLER_97_369 ();
 FILLCELL_X4 FILLER_97_412 ();
 FILLCELL_X16 FILLER_97_433 ();
 FILLCELL_X1 FILLER_97_449 ();
 FILLCELL_X32 FILLER_97_457 ();
 FILLCELL_X8 FILLER_97_489 ();
 FILLCELL_X4 FILLER_97_497 ();
 FILLCELL_X1 FILLER_97_501 ();
 FILLCELL_X2 FILLER_97_506 ();
 FILLCELL_X1 FILLER_97_508 ();
 FILLCELL_X2 FILLER_97_516 ();
 FILLCELL_X1 FILLER_97_532 ();
 FILLCELL_X1 FILLER_97_543 ();
 FILLCELL_X4 FILLER_97_559 ();
 FILLCELL_X16 FILLER_97_573 ();
 FILLCELL_X8 FILLER_97_589 ();
 FILLCELL_X4 FILLER_97_597 ();
 FILLCELL_X2 FILLER_97_601 ();
 FILLCELL_X16 FILLER_97_607 ();
 FILLCELL_X8 FILLER_97_623 ();
 FILLCELL_X2 FILLER_97_631 ();
 FILLCELL_X1 FILLER_97_633 ();
 FILLCELL_X2 FILLER_97_655 ();
 FILLCELL_X4 FILLER_97_672 ();
 FILLCELL_X1 FILLER_97_676 ();
 FILLCELL_X1 FILLER_97_679 ();
 FILLCELL_X8 FILLER_97_712 ();
 FILLCELL_X4 FILLER_97_720 ();
 FILLCELL_X2 FILLER_97_724 ();
 FILLCELL_X1 FILLER_97_726 ();
 FILLCELL_X4 FILLER_97_737 ();
 FILLCELL_X2 FILLER_97_741 ();
 FILLCELL_X4 FILLER_97_774 ();
 FILLCELL_X2 FILLER_97_778 ();
 FILLCELL_X1 FILLER_97_780 ();
 FILLCELL_X4 FILLER_97_788 ();
 FILLCELL_X8 FILLER_97_795 ();
 FILLCELL_X4 FILLER_97_803 ();
 FILLCELL_X2 FILLER_97_807 ();
 FILLCELL_X2 FILLER_97_816 ();
 FILLCELL_X8 FILLER_97_848 ();
 FILLCELL_X2 FILLER_97_856 ();
 FILLCELL_X1 FILLER_97_858 ();
 FILLCELL_X1 FILLER_97_863 ();
 FILLCELL_X4 FILLER_97_879 ();
 FILLCELL_X1 FILLER_97_885 ();
 FILLCELL_X2 FILLER_97_898 ();
 FILLCELL_X2 FILLER_97_920 ();
 FILLCELL_X2 FILLER_97_926 ();
 FILLCELL_X1 FILLER_97_928 ();
 FILLCELL_X1 FILLER_97_933 ();
 FILLCELL_X8 FILLER_97_959 ();
 FILLCELL_X4 FILLER_97_974 ();
 FILLCELL_X1 FILLER_97_978 ();
 FILLCELL_X8 FILLER_97_993 ();
 FILLCELL_X4 FILLER_97_1001 ();
 FILLCELL_X2 FILLER_97_1005 ();
 FILLCELL_X16 FILLER_97_1014 ();
 FILLCELL_X2 FILLER_97_1030 ();
 FILLCELL_X8 FILLER_97_1039 ();
 FILLCELL_X4 FILLER_97_1061 ();
 FILLCELL_X1 FILLER_97_1065 ();
 FILLCELL_X2 FILLER_97_1083 ();
 FILLCELL_X2 FILLER_97_1089 ();
 FILLCELL_X1 FILLER_97_1091 ();
 FILLCELL_X1 FILLER_97_1096 ();
 FILLCELL_X8 FILLER_97_1117 ();
 FILLCELL_X4 FILLER_97_1125 ();
 FILLCELL_X2 FILLER_97_1129 ();
 FILLCELL_X2 FILLER_97_1148 ();
 FILLCELL_X1 FILLER_97_1150 ();
 FILLCELL_X8 FILLER_97_1156 ();
 FILLCELL_X4 FILLER_97_1164 ();
 FILLCELL_X1 FILLER_97_1168 ();
 FILLCELL_X4 FILLER_97_1188 ();
 FILLCELL_X1 FILLER_97_1192 ();
 FILLCELL_X8 FILLER_97_1199 ();
 FILLCELL_X2 FILLER_97_1207 ();
 FILLCELL_X32 FILLER_98_1 ();
 FILLCELL_X32 FILLER_98_36 ();
 FILLCELL_X32 FILLER_98_68 ();
 FILLCELL_X8 FILLER_98_100 ();
 FILLCELL_X4 FILLER_98_108 ();
 FILLCELL_X2 FILLER_98_112 ();
 FILLCELL_X1 FILLER_98_114 ();
 FILLCELL_X8 FILLER_98_139 ();
 FILLCELL_X1 FILLER_98_147 ();
 FILLCELL_X1 FILLER_98_177 ();
 FILLCELL_X4 FILLER_98_194 ();
 FILLCELL_X2 FILLER_98_198 ();
 FILLCELL_X4 FILLER_98_219 ();
 FILLCELL_X4 FILLER_98_234 ();
 FILLCELL_X2 FILLER_98_247 ();
 FILLCELL_X1 FILLER_98_249 ();
 FILLCELL_X4 FILLER_98_257 ();
 FILLCELL_X2 FILLER_98_261 ();
 FILLCELL_X1 FILLER_98_263 ();
 FILLCELL_X16 FILLER_98_273 ();
 FILLCELL_X4 FILLER_98_289 ();
 FILLCELL_X1 FILLER_98_293 ();
 FILLCELL_X8 FILLER_98_301 ();
 FILLCELL_X4 FILLER_98_309 ();
 FILLCELL_X1 FILLER_98_313 ();
 FILLCELL_X4 FILLER_98_333 ();
 FILLCELL_X2 FILLER_98_358 ();
 FILLCELL_X1 FILLER_98_360 ();
 FILLCELL_X1 FILLER_98_370 ();
 FILLCELL_X4 FILLER_98_396 ();
 FILLCELL_X1 FILLER_98_400 ();
 FILLCELL_X16 FILLER_98_423 ();
 FILLCELL_X4 FILLER_98_439 ();
 FILLCELL_X32 FILLER_98_448 ();
 FILLCELL_X16 FILLER_98_480 ();
 FILLCELL_X8 FILLER_98_496 ();
 FILLCELL_X4 FILLER_98_504 ();
 FILLCELL_X2 FILLER_98_508 ();
 FILLCELL_X2 FILLER_98_514 ();
 FILLCELL_X1 FILLER_98_516 ();
 FILLCELL_X8 FILLER_98_523 ();
 FILLCELL_X4 FILLER_98_531 ();
 FILLCELL_X1 FILLER_98_535 ();
 FILLCELL_X2 FILLER_98_547 ();
 FILLCELL_X1 FILLER_98_549 ();
 FILLCELL_X8 FILLER_98_559 ();
 FILLCELL_X4 FILLER_98_567 ();
 FILLCELL_X2 FILLER_98_571 ();
 FILLCELL_X1 FILLER_98_573 ();
 FILLCELL_X8 FILLER_98_581 ();
 FILLCELL_X2 FILLER_98_589 ();
 FILLCELL_X4 FILLER_98_598 ();
 FILLCELL_X1 FILLER_98_613 ();
 FILLCELL_X2 FILLER_98_632 ();
 FILLCELL_X4 FILLER_98_647 ();
 FILLCELL_X8 FILLER_98_698 ();
 FILLCELL_X4 FILLER_98_706 ();
 FILLCELL_X4 FILLER_98_713 ();
 FILLCELL_X2 FILLER_98_717 ();
 FILLCELL_X8 FILLER_98_753 ();
 FILLCELL_X2 FILLER_98_761 ();
 FILLCELL_X4 FILLER_98_769 ();
 FILLCELL_X1 FILLER_98_773 ();
 FILLCELL_X8 FILLER_98_793 ();
 FILLCELL_X4 FILLER_98_801 ();
 FILLCELL_X2 FILLER_98_838 ();
 FILLCELL_X1 FILLER_98_845 ();
 FILLCELL_X8 FILLER_98_870 ();
 FILLCELL_X4 FILLER_98_878 ();
 FILLCELL_X2 FILLER_98_882 ();
 FILLCELL_X1 FILLER_98_884 ();
 FILLCELL_X1 FILLER_98_902 ();
 FILLCELL_X2 FILLER_98_912 ();
 FILLCELL_X1 FILLER_98_914 ();
 FILLCELL_X2 FILLER_98_934 ();
 FILLCELL_X1 FILLER_98_945 ();
 FILLCELL_X4 FILLER_98_954 ();
 FILLCELL_X2 FILLER_98_958 ();
 FILLCELL_X1 FILLER_98_960 ();
 FILLCELL_X8 FILLER_98_990 ();
 FILLCELL_X1 FILLER_98_1011 ();
 FILLCELL_X1 FILLER_98_1026 ();
 FILLCELL_X2 FILLER_98_1047 ();
 FILLCELL_X2 FILLER_98_1059 ();
 FILLCELL_X4 FILLER_98_1103 ();
 FILLCELL_X1 FILLER_98_1107 ();
 FILLCELL_X4 FILLER_98_1116 ();
 FILLCELL_X2 FILLER_98_1120 ();
 FILLCELL_X2 FILLER_98_1139 ();
 FILLCELL_X1 FILLER_98_1150 ();
 FILLCELL_X8 FILLER_98_1154 ();
 FILLCELL_X2 FILLER_98_1169 ();
 FILLCELL_X1 FILLER_98_1171 ();
 FILLCELL_X8 FILLER_98_1196 ();
 FILLCELL_X4 FILLER_98_1204 ();
 FILLCELL_X1 FILLER_98_1208 ();
 FILLCELL_X32 FILLER_99_1 ();
 FILLCELL_X32 FILLER_99_33 ();
 FILLCELL_X32 FILLER_99_65 ();
 FILLCELL_X16 FILLER_99_97 ();
 FILLCELL_X1 FILLER_99_147 ();
 FILLCELL_X2 FILLER_99_165 ();
 FILLCELL_X1 FILLER_99_203 ();
 FILLCELL_X8 FILLER_99_215 ();
 FILLCELL_X4 FILLER_99_223 ();
 FILLCELL_X16 FILLER_99_232 ();
 FILLCELL_X2 FILLER_99_248 ();
 FILLCELL_X2 FILLER_99_263 ();
 FILLCELL_X1 FILLER_99_265 ();
 FILLCELL_X1 FILLER_99_295 ();
 FILLCELL_X8 FILLER_99_322 ();
 FILLCELL_X4 FILLER_99_330 ();
 FILLCELL_X1 FILLER_99_334 ();
 FILLCELL_X2 FILLER_99_352 ();
 FILLCELL_X4 FILLER_99_361 ();
 FILLCELL_X1 FILLER_99_365 ();
 FILLCELL_X8 FILLER_99_374 ();
 FILLCELL_X4 FILLER_99_385 ();
 FILLCELL_X8 FILLER_99_416 ();
 FILLCELL_X4 FILLER_99_424 ();
 FILLCELL_X2 FILLER_99_428 ();
 FILLCELL_X16 FILLER_99_447 ();
 FILLCELL_X8 FILLER_99_463 ();
 FILLCELL_X4 FILLER_99_471 ();
 FILLCELL_X1 FILLER_99_475 ();
 FILLCELL_X8 FILLER_99_493 ();
 FILLCELL_X4 FILLER_99_501 ();
 FILLCELL_X16 FILLER_99_513 ();
 FILLCELL_X1 FILLER_99_529 ();
 FILLCELL_X8 FILLER_99_543 ();
 FILLCELL_X2 FILLER_99_551 ();
 FILLCELL_X8 FILLER_99_559 ();
 FILLCELL_X1 FILLER_99_567 ();
 FILLCELL_X4 FILLER_99_596 ();
 FILLCELL_X1 FILLER_99_611 ();
 FILLCELL_X4 FILLER_99_616 ();
 FILLCELL_X2 FILLER_99_620 ();
 FILLCELL_X1 FILLER_99_622 ();
 FILLCELL_X2 FILLER_99_634 ();
 FILLCELL_X1 FILLER_99_640 ();
 FILLCELL_X2 FILLER_99_656 ();
 FILLCELL_X1 FILLER_99_658 ();
 FILLCELL_X2 FILLER_99_666 ();
 FILLCELL_X1 FILLER_99_668 ();
 FILLCELL_X8 FILLER_99_697 ();
 FILLCELL_X1 FILLER_99_705 ();
 FILLCELL_X4 FILLER_99_720 ();
 FILLCELL_X1 FILLER_99_724 ();
 FILLCELL_X4 FILLER_99_728 ();
 FILLCELL_X4 FILLER_99_756 ();
 FILLCELL_X2 FILLER_99_780 ();
 FILLCELL_X1 FILLER_99_782 ();
 FILLCELL_X16 FILLER_99_800 ();
 FILLCELL_X2 FILLER_99_816 ();
 FILLCELL_X1 FILLER_99_843 ();
 FILLCELL_X1 FILLER_99_850 ();
 FILLCELL_X1 FILLER_99_870 ();
 FILLCELL_X16 FILLER_99_879 ();
 FILLCELL_X2 FILLER_99_895 ();
 FILLCELL_X4 FILLER_99_907 ();
 FILLCELL_X1 FILLER_99_915 ();
 FILLCELL_X2 FILLER_99_919 ();
 FILLCELL_X2 FILLER_99_930 ();
 FILLCELL_X1 FILLER_99_932 ();
 FILLCELL_X8 FILLER_99_981 ();
 FILLCELL_X4 FILLER_99_989 ();
 FILLCELL_X2 FILLER_99_993 ();
 FILLCELL_X16 FILLER_99_1017 ();
 FILLCELL_X4 FILLER_99_1033 ();
 FILLCELL_X1 FILLER_99_1037 ();
 FILLCELL_X2 FILLER_99_1061 ();
 FILLCELL_X1 FILLER_99_1076 ();
 FILLCELL_X4 FILLER_99_1088 ();
 FILLCELL_X2 FILLER_99_1096 ();
 FILLCELL_X1 FILLER_99_1098 ();
 FILLCELL_X1 FILLER_99_1108 ();
 FILLCELL_X4 FILLER_99_1172 ();
 FILLCELL_X2 FILLER_99_1176 ();
 FILLCELL_X2 FILLER_99_1195 ();
 FILLCELL_X1 FILLER_99_1197 ();
 FILLCELL_X2 FILLER_99_1204 ();
 FILLCELL_X32 FILLER_100_1 ();
 FILLCELL_X32 FILLER_100_33 ();
 FILLCELL_X16 FILLER_100_65 ();
 FILLCELL_X1 FILLER_100_81 ();
 FILLCELL_X16 FILLER_100_99 ();
 FILLCELL_X1 FILLER_100_115 ();
 FILLCELL_X4 FILLER_100_123 ();
 FILLCELL_X1 FILLER_100_134 ();
 FILLCELL_X4 FILLER_100_148 ();
 FILLCELL_X2 FILLER_100_163 ();
 FILLCELL_X2 FILLER_100_187 ();
 FILLCELL_X1 FILLER_100_215 ();
 FILLCELL_X2 FILLER_100_226 ();
 FILLCELL_X32 FILLER_100_243 ();
 FILLCELL_X2 FILLER_100_275 ();
 FILLCELL_X1 FILLER_100_277 ();
 FILLCELL_X2 FILLER_100_296 ();
 FILLCELL_X1 FILLER_100_298 ();
 FILLCELL_X8 FILLER_100_301 ();
 FILLCELL_X2 FILLER_100_309 ();
 FILLCELL_X2 FILLER_100_328 ();
 FILLCELL_X1 FILLER_100_330 ();
 FILLCELL_X2 FILLER_100_362 ();
 FILLCELL_X8 FILLER_100_393 ();
 FILLCELL_X1 FILLER_100_401 ();
 FILLCELL_X1 FILLER_100_423 ();
 FILLCELL_X32 FILLER_100_467 ();
 FILLCELL_X2 FILLER_100_499 ();
 FILLCELL_X4 FILLER_100_507 ();
 FILLCELL_X2 FILLER_100_511 ();
 FILLCELL_X1 FILLER_100_513 ();
 FILLCELL_X1 FILLER_100_519 ();
 FILLCELL_X16 FILLER_100_530 ();
 FILLCELL_X8 FILLER_100_546 ();
 FILLCELL_X2 FILLER_100_554 ();
 FILLCELL_X4 FILLER_100_559 ();
 FILLCELL_X4 FILLER_100_566 ();
 FILLCELL_X2 FILLER_100_570 ();
 FILLCELL_X1 FILLER_100_572 ();
 FILLCELL_X2 FILLER_100_602 ();
 FILLCELL_X8 FILLER_100_615 ();
 FILLCELL_X2 FILLER_100_623 ();
 FILLCELL_X1 FILLER_100_625 ();
 FILLCELL_X1 FILLER_100_630 ();
 FILLCELL_X4 FILLER_100_632 ();
 FILLCELL_X1 FILLER_100_648 ();
 FILLCELL_X4 FILLER_100_656 ();
 FILLCELL_X1 FILLER_100_660 ();
 FILLCELL_X1 FILLER_100_689 ();
 FILLCELL_X2 FILLER_100_702 ();
 FILLCELL_X1 FILLER_100_704 ();
 FILLCELL_X1 FILLER_100_724 ();
 FILLCELL_X4 FILLER_100_733 ();
 FILLCELL_X2 FILLER_100_737 ();
 FILLCELL_X4 FILLER_100_743 ();
 FILLCELL_X2 FILLER_100_747 ();
 FILLCELL_X2 FILLER_100_755 ();
 FILLCELL_X4 FILLER_100_775 ();
 FILLCELL_X4 FILLER_100_786 ();
 FILLCELL_X1 FILLER_100_797 ();
 FILLCELL_X4 FILLER_100_815 ();
 FILLCELL_X2 FILLER_100_819 ();
 FILLCELL_X1 FILLER_100_821 ();
 FILLCELL_X2 FILLER_100_839 ();
 FILLCELL_X1 FILLER_100_858 ();
 FILLCELL_X8 FILLER_100_884 ();
 FILLCELL_X2 FILLER_100_892 ();
 FILLCELL_X4 FILLER_100_920 ();
 FILLCELL_X1 FILLER_100_924 ();
 FILLCELL_X4 FILLER_100_939 ();
 FILLCELL_X8 FILLER_100_956 ();
 FILLCELL_X8 FILLER_100_978 ();
 FILLCELL_X1 FILLER_100_986 ();
 FILLCELL_X2 FILLER_100_1000 ();
 FILLCELL_X1 FILLER_100_1002 ();
 FILLCELL_X1 FILLER_100_1020 ();
 FILLCELL_X1 FILLER_100_1068 ();
 FILLCELL_X1 FILLER_100_1104 ();
 FILLCELL_X8 FILLER_100_1109 ();
 FILLCELL_X2 FILLER_100_1130 ();
 FILLCELL_X1 FILLER_100_1136 ();
 FILLCELL_X4 FILLER_100_1155 ();
 FILLCELL_X2 FILLER_100_1159 ();
 FILLCELL_X1 FILLER_100_1161 ();
 FILLCELL_X1 FILLER_100_1175 ();
 FILLCELL_X8 FILLER_100_1184 ();
 FILLCELL_X1 FILLER_100_1192 ();
 FILLCELL_X8 FILLER_100_1197 ();
 FILLCELL_X4 FILLER_100_1205 ();
 FILLCELL_X16 FILLER_101_1 ();
 FILLCELL_X4 FILLER_101_17 ();
 FILLCELL_X32 FILLER_101_24 ();
 FILLCELL_X32 FILLER_101_56 ();
 FILLCELL_X16 FILLER_101_88 ();
 FILLCELL_X4 FILLER_101_104 ();
 FILLCELL_X1 FILLER_101_108 ();
 FILLCELL_X1 FILLER_101_129 ();
 FILLCELL_X1 FILLER_101_142 ();
 FILLCELL_X1 FILLER_101_150 ();
 FILLCELL_X2 FILLER_101_164 ();
 FILLCELL_X2 FILLER_101_171 ();
 FILLCELL_X1 FILLER_101_173 ();
 FILLCELL_X1 FILLER_101_180 ();
 FILLCELL_X2 FILLER_101_223 ();
 FILLCELL_X1 FILLER_101_230 ();
 FILLCELL_X8 FILLER_101_263 ();
 FILLCELL_X2 FILLER_101_271 ();
 FILLCELL_X1 FILLER_101_273 ();
 FILLCELL_X8 FILLER_101_283 ();
 FILLCELL_X1 FILLER_101_291 ();
 FILLCELL_X8 FILLER_101_305 ();
 FILLCELL_X2 FILLER_101_313 ();
 FILLCELL_X1 FILLER_101_315 ();
 FILLCELL_X2 FILLER_101_354 ();
 FILLCELL_X1 FILLER_101_356 ();
 FILLCELL_X2 FILLER_101_364 ();
 FILLCELL_X1 FILLER_101_366 ();
 FILLCELL_X1 FILLER_101_370 ();
 FILLCELL_X4 FILLER_101_384 ();
 FILLCELL_X1 FILLER_101_407 ();
 FILLCELL_X1 FILLER_101_411 ();
 FILLCELL_X4 FILLER_101_437 ();
 FILLCELL_X2 FILLER_101_441 ();
 FILLCELL_X1 FILLER_101_443 ();
 FILLCELL_X16 FILLER_101_466 ();
 FILLCELL_X1 FILLER_101_482 ();
 FILLCELL_X16 FILLER_101_487 ();
 FILLCELL_X2 FILLER_101_503 ();
 FILLCELL_X1 FILLER_101_505 ();
 FILLCELL_X1 FILLER_101_524 ();
 FILLCELL_X4 FILLER_101_534 ();
 FILLCELL_X2 FILLER_101_538 ();
 FILLCELL_X8 FILLER_101_544 ();
 FILLCELL_X4 FILLER_101_552 ();
 FILLCELL_X32 FILLER_101_560 ();
 FILLCELL_X16 FILLER_101_592 ();
 FILLCELL_X8 FILLER_101_608 ();
 FILLCELL_X4 FILLER_101_616 ();
 FILLCELL_X2 FILLER_101_620 ();
 FILLCELL_X1 FILLER_101_622 ();
 FILLCELL_X1 FILLER_101_639 ();
 FILLCELL_X8 FILLER_101_655 ();
 FILLCELL_X2 FILLER_101_663 ();
 FILLCELL_X1 FILLER_101_665 ();
 FILLCELL_X4 FILLER_101_677 ();
 FILLCELL_X16 FILLER_101_692 ();
 FILLCELL_X8 FILLER_101_708 ();
 FILLCELL_X1 FILLER_101_716 ();
 FILLCELL_X1 FILLER_101_722 ();
 FILLCELL_X8 FILLER_101_737 ();
 FILLCELL_X2 FILLER_101_745 ();
 FILLCELL_X4 FILLER_101_769 ();
 FILLCELL_X1 FILLER_101_773 ();
 FILLCELL_X16 FILLER_101_808 ();
 FILLCELL_X8 FILLER_101_824 ();
 FILLCELL_X4 FILLER_101_832 ();
 FILLCELL_X8 FILLER_101_888 ();
 FILLCELL_X4 FILLER_101_918 ();
 FILLCELL_X2 FILLER_101_922 ();
 FILLCELL_X1 FILLER_101_924 ();
 FILLCELL_X1 FILLER_101_936 ();
 FILLCELL_X1 FILLER_101_941 ();
 FILLCELL_X32 FILLER_101_945 ();
 FILLCELL_X1 FILLER_101_977 ();
 FILLCELL_X8 FILLER_101_991 ();
 FILLCELL_X4 FILLER_101_999 ();
 FILLCELL_X1 FILLER_101_1017 ();
 FILLCELL_X4 FILLER_101_1040 ();
 FILLCELL_X2 FILLER_101_1044 ();
 FILLCELL_X2 FILLER_101_1063 ();
 FILLCELL_X2 FILLER_101_1081 ();
 FILLCELL_X2 FILLER_101_1092 ();
 FILLCELL_X1 FILLER_101_1094 ();
 FILLCELL_X2 FILLER_101_1172 ();
 FILLCELL_X2 FILLER_101_1178 ();
 FILLCELL_X2 FILLER_101_1191 ();
 FILLCELL_X4 FILLER_101_1196 ();
 FILLCELL_X4 FILLER_101_1203 ();
 FILLCELL_X2 FILLER_101_1207 ();
 FILLCELL_X32 FILLER_102_1 ();
 FILLCELL_X32 FILLER_102_33 ();
 FILLCELL_X32 FILLER_102_65 ();
 FILLCELL_X2 FILLER_102_97 ();
 FILLCELL_X1 FILLER_102_99 ();
 FILLCELL_X4 FILLER_102_107 ();
 FILLCELL_X1 FILLER_102_111 ();
 FILLCELL_X4 FILLER_102_125 ();
 FILLCELL_X2 FILLER_102_129 ();
 FILLCELL_X4 FILLER_102_155 ();
 FILLCELL_X4 FILLER_102_163 ();
 FILLCELL_X2 FILLER_102_173 ();
 FILLCELL_X1 FILLER_102_175 ();
 FILLCELL_X1 FILLER_102_189 ();
 FILLCELL_X2 FILLER_102_196 ();
 FILLCELL_X1 FILLER_102_198 ();
 FILLCELL_X1 FILLER_102_231 ();
 FILLCELL_X1 FILLER_102_248 ();
 FILLCELL_X2 FILLER_102_261 ();
 FILLCELL_X4 FILLER_102_270 ();
 FILLCELL_X16 FILLER_102_283 ();
 FILLCELL_X4 FILLER_102_304 ();
 FILLCELL_X1 FILLER_102_308 ();
 FILLCELL_X1 FILLER_102_325 ();
 FILLCELL_X1 FILLER_102_335 ();
 FILLCELL_X1 FILLER_102_339 ();
 FILLCELL_X2 FILLER_102_343 ();
 FILLCELL_X1 FILLER_102_348 ();
 FILLCELL_X4 FILLER_102_351 ();
 FILLCELL_X4 FILLER_102_372 ();
 FILLCELL_X1 FILLER_102_376 ();
 FILLCELL_X8 FILLER_102_431 ();
 FILLCELL_X4 FILLER_102_439 ();
 FILLCELL_X32 FILLER_102_447 ();
 FILLCELL_X16 FILLER_102_479 ();
 FILLCELL_X4 FILLER_102_495 ();
 FILLCELL_X2 FILLER_102_499 ();
 FILLCELL_X1 FILLER_102_505 ();
 FILLCELL_X2 FILLER_102_509 ();
 FILLCELL_X1 FILLER_102_514 ();
 FILLCELL_X8 FILLER_102_523 ();
 FILLCELL_X4 FILLER_102_531 ();
 FILLCELL_X1 FILLER_102_539 ();
 FILLCELL_X1 FILLER_102_551 ();
 FILLCELL_X1 FILLER_102_555 ();
 FILLCELL_X8 FILLER_102_567 ();
 FILLCELL_X2 FILLER_102_575 ();
 FILLCELL_X8 FILLER_102_582 ();
 FILLCELL_X2 FILLER_102_590 ();
 FILLCELL_X16 FILLER_102_596 ();
 FILLCELL_X4 FILLER_102_612 ();
 FILLCELL_X2 FILLER_102_616 ();
 FILLCELL_X1 FILLER_102_618 ();
 FILLCELL_X4 FILLER_102_627 ();
 FILLCELL_X1 FILLER_102_632 ();
 FILLCELL_X8 FILLER_102_644 ();
 FILLCELL_X2 FILLER_102_652 ();
 FILLCELL_X16 FILLER_102_658 ();
 FILLCELL_X2 FILLER_102_674 ();
 FILLCELL_X2 FILLER_102_680 ();
 FILLCELL_X1 FILLER_102_682 ();
 FILLCELL_X16 FILLER_102_687 ();
 FILLCELL_X8 FILLER_102_703 ();
 FILLCELL_X4 FILLER_102_711 ();
 FILLCELL_X1 FILLER_102_715 ();
 FILLCELL_X4 FILLER_102_719 ();
 FILLCELL_X2 FILLER_102_723 ();
 FILLCELL_X4 FILLER_102_736 ();
 FILLCELL_X1 FILLER_102_740 ();
 FILLCELL_X1 FILLER_102_744 ();
 FILLCELL_X1 FILLER_102_776 ();
 FILLCELL_X8 FILLER_102_783 ();
 FILLCELL_X1 FILLER_102_791 ();
 FILLCELL_X16 FILLER_102_795 ();
 FILLCELL_X2 FILLER_102_811 ();
 FILLCELL_X4 FILLER_102_842 ();
 FILLCELL_X2 FILLER_102_846 ();
 FILLCELL_X1 FILLER_102_848 ();
 FILLCELL_X4 FILLER_102_856 ();
 FILLCELL_X1 FILLER_102_860 ();
 FILLCELL_X8 FILLER_102_883 ();
 FILLCELL_X2 FILLER_102_891 ();
 FILLCELL_X2 FILLER_102_905 ();
 FILLCELL_X1 FILLER_102_926 ();
 FILLCELL_X1 FILLER_102_947 ();
 FILLCELL_X4 FILLER_102_951 ();
 FILLCELL_X1 FILLER_102_955 ();
 FILLCELL_X1 FILLER_102_962 ();
 FILLCELL_X4 FILLER_102_985 ();
 FILLCELL_X2 FILLER_102_1015 ();
 FILLCELL_X2 FILLER_102_1031 ();
 FILLCELL_X2 FILLER_102_1036 ();
 FILLCELL_X4 FILLER_102_1049 ();
 FILLCELL_X4 FILLER_102_1056 ();
 FILLCELL_X2 FILLER_102_1070 ();
 FILLCELL_X16 FILLER_102_1088 ();
 FILLCELL_X1 FILLER_102_1104 ();
 FILLCELL_X4 FILLER_102_1110 ();
 FILLCELL_X2 FILLER_102_1114 ();
 FILLCELL_X1 FILLER_102_1116 ();
 FILLCELL_X1 FILLER_102_1130 ();
 FILLCELL_X1 FILLER_102_1142 ();
 FILLCELL_X2 FILLER_102_1163 ();
 FILLCELL_X1 FILLER_102_1185 ();
 FILLCELL_X16 FILLER_102_1193 ();
 FILLCELL_X16 FILLER_103_1 ();
 FILLCELL_X8 FILLER_103_17 ();
 FILLCELL_X32 FILLER_103_28 ();
 FILLCELL_X32 FILLER_103_60 ();
 FILLCELL_X8 FILLER_103_92 ();
 FILLCELL_X2 FILLER_103_100 ();
 FILLCELL_X1 FILLER_103_102 ();
 FILLCELL_X1 FILLER_103_110 ();
 FILLCELL_X1 FILLER_103_118 ();
 FILLCELL_X1 FILLER_103_127 ();
 FILLCELL_X2 FILLER_103_132 ();
 FILLCELL_X2 FILLER_103_161 ();
 FILLCELL_X2 FILLER_103_166 ();
 FILLCELL_X4 FILLER_103_173 ();
 FILLCELL_X2 FILLER_103_177 ();
 FILLCELL_X4 FILLER_103_188 ();
 FILLCELL_X2 FILLER_103_192 ();
 FILLCELL_X1 FILLER_103_200 ();
 FILLCELL_X1 FILLER_103_220 ();
 FILLCELL_X1 FILLER_103_225 ();
 FILLCELL_X1 FILLER_103_236 ();
 FILLCELL_X2 FILLER_103_259 ();
 FILLCELL_X32 FILLER_103_282 ();
 FILLCELL_X2 FILLER_103_314 ();
 FILLCELL_X4 FILLER_103_328 ();
 FILLCELL_X1 FILLER_103_332 ();
 FILLCELL_X16 FILLER_103_350 ();
 FILLCELL_X8 FILLER_103_366 ();
 FILLCELL_X1 FILLER_103_374 ();
 FILLCELL_X1 FILLER_103_393 ();
 FILLCELL_X1 FILLER_103_420 ();
 FILLCELL_X8 FILLER_103_425 ();
 FILLCELL_X1 FILLER_103_433 ();
 FILLCELL_X32 FILLER_103_451 ();
 FILLCELL_X16 FILLER_103_483 ();
 FILLCELL_X4 FILLER_103_499 ();
 FILLCELL_X2 FILLER_103_503 ();
 FILLCELL_X1 FILLER_103_505 ();
 FILLCELL_X2 FILLER_103_537 ();
 FILLCELL_X2 FILLER_103_543 ();
 FILLCELL_X16 FILLER_103_559 ();
 FILLCELL_X2 FILLER_103_579 ();
 FILLCELL_X1 FILLER_103_581 ();
 FILLCELL_X1 FILLER_103_589 ();
 FILLCELL_X16 FILLER_103_600 ();
 FILLCELL_X8 FILLER_103_616 ();
 FILLCELL_X8 FILLER_103_628 ();
 FILLCELL_X4 FILLER_103_636 ();
 FILLCELL_X2 FILLER_103_640 ();
 FILLCELL_X1 FILLER_103_642 ();
 FILLCELL_X8 FILLER_103_648 ();
 FILLCELL_X1 FILLER_103_656 ();
 FILLCELL_X8 FILLER_103_661 ();
 FILLCELL_X1 FILLER_103_669 ();
 FILLCELL_X16 FILLER_103_691 ();
 FILLCELL_X4 FILLER_103_707 ();
 FILLCELL_X2 FILLER_103_711 ();
 FILLCELL_X16 FILLER_103_730 ();
 FILLCELL_X8 FILLER_103_750 ();
 FILLCELL_X2 FILLER_103_758 ();
 FILLCELL_X1 FILLER_103_760 ();
 FILLCELL_X16 FILLER_103_805 ();
 FILLCELL_X4 FILLER_103_821 ();
 FILLCELL_X2 FILLER_103_847 ();
 FILLCELL_X1 FILLER_103_859 ();
 FILLCELL_X8 FILLER_103_869 ();
 FILLCELL_X2 FILLER_103_877 ();
 FILLCELL_X16 FILLER_103_892 ();
 FILLCELL_X8 FILLER_103_908 ();
 FILLCELL_X4 FILLER_103_916 ();
 FILLCELL_X1 FILLER_103_920 ();
 FILLCELL_X4 FILLER_103_928 ();
 FILLCELL_X8 FILLER_103_945 ();
 FILLCELL_X2 FILLER_103_953 ();
 FILLCELL_X1 FILLER_103_955 ();
 FILLCELL_X2 FILLER_103_959 ();
 FILLCELL_X1 FILLER_103_961 ();
 FILLCELL_X16 FILLER_103_969 ();
 FILLCELL_X4 FILLER_103_985 ();
 FILLCELL_X2 FILLER_103_1001 ();
 FILLCELL_X1 FILLER_103_1003 ();
 FILLCELL_X1 FILLER_103_1031 ();
 FILLCELL_X8 FILLER_103_1036 ();
 FILLCELL_X2 FILLER_103_1044 ();
 FILLCELL_X1 FILLER_103_1046 ();
 FILLCELL_X4 FILLER_103_1051 ();
 FILLCELL_X2 FILLER_103_1055 ();
 FILLCELL_X1 FILLER_103_1061 ();
 FILLCELL_X2 FILLER_103_1065 ();
 FILLCELL_X8 FILLER_103_1070 ();
 FILLCELL_X4 FILLER_103_1078 ();
 FILLCELL_X16 FILLER_103_1093 ();
 FILLCELL_X8 FILLER_103_1116 ();
 FILLCELL_X1 FILLER_103_1124 ();
 FILLCELL_X1 FILLER_103_1137 ();
 FILLCELL_X8 FILLER_103_1185 ();
 FILLCELL_X4 FILLER_103_1193 ();
 FILLCELL_X8 FILLER_103_1200 ();
 FILLCELL_X1 FILLER_103_1208 ();
 FILLCELL_X32 FILLER_104_1 ();
 FILLCELL_X32 FILLER_104_33 ();
 FILLCELL_X32 FILLER_104_65 ();
 FILLCELL_X8 FILLER_104_97 ();
 FILLCELL_X4 FILLER_104_105 ();
 FILLCELL_X1 FILLER_104_109 ();
 FILLCELL_X2 FILLER_104_115 ();
 FILLCELL_X4 FILLER_104_121 ();
 FILLCELL_X2 FILLER_104_125 ();
 FILLCELL_X2 FILLER_104_140 ();
 FILLCELL_X2 FILLER_104_158 ();
 FILLCELL_X1 FILLER_104_160 ();
 FILLCELL_X4 FILLER_104_165 ();
 FILLCELL_X2 FILLER_104_169 ();
 FILLCELL_X1 FILLER_104_186 ();
 FILLCELL_X1 FILLER_104_198 ();
 FILLCELL_X1 FILLER_104_203 ();
 FILLCELL_X1 FILLER_104_209 ();
 FILLCELL_X2 FILLER_104_230 ();
 FILLCELL_X1 FILLER_104_232 ();
 FILLCELL_X2 FILLER_104_235 ();
 FILLCELL_X2 FILLER_104_265 ();
 FILLCELL_X1 FILLER_104_267 ();
 FILLCELL_X16 FILLER_104_322 ();
 FILLCELL_X2 FILLER_104_338 ();
 FILLCELL_X1 FILLER_104_340 ();
 FILLCELL_X16 FILLER_104_352 ();
 FILLCELL_X8 FILLER_104_368 ();
 FILLCELL_X1 FILLER_104_376 ();
 FILLCELL_X4 FILLER_104_394 ();
 FILLCELL_X1 FILLER_104_398 ();
 FILLCELL_X2 FILLER_104_411 ();
 FILLCELL_X2 FILLER_104_418 ();
 FILLCELL_X2 FILLER_104_433 ();
 FILLCELL_X8 FILLER_104_451 ();
 FILLCELL_X4 FILLER_104_459 ();
 FILLCELL_X2 FILLER_104_463 ();
 FILLCELL_X1 FILLER_104_465 ();
 FILLCELL_X8 FILLER_104_471 ();
 FILLCELL_X4 FILLER_104_479 ();
 FILLCELL_X1 FILLER_104_483 ();
 FILLCELL_X4 FILLER_104_501 ();
 FILLCELL_X2 FILLER_104_518 ();
 FILLCELL_X2 FILLER_104_558 ();
 FILLCELL_X4 FILLER_104_570 ();
 FILLCELL_X2 FILLER_104_585 ();
 FILLCELL_X1 FILLER_104_587 ();
 FILLCELL_X2 FILLER_104_599 ();
 FILLCELL_X1 FILLER_104_601 ();
 FILLCELL_X4 FILLER_104_616 ();
 FILLCELL_X2 FILLER_104_620 ();
 FILLCELL_X4 FILLER_104_626 ();
 FILLCELL_X1 FILLER_104_630 ();
 FILLCELL_X8 FILLER_104_632 ();
 FILLCELL_X2 FILLER_104_644 ();
 FILLCELL_X1 FILLER_104_646 ();
 FILLCELL_X2 FILLER_104_670 ();
 FILLCELL_X1 FILLER_104_672 ();
 FILLCELL_X16 FILLER_104_699 ();
 FILLCELL_X4 FILLER_104_715 ();
 FILLCELL_X2 FILLER_104_719 ();
 FILLCELL_X8 FILLER_104_760 ();
 FILLCELL_X16 FILLER_104_784 ();
 FILLCELL_X4 FILLER_104_800 ();
 FILLCELL_X2 FILLER_104_804 ();
 FILLCELL_X16 FILLER_104_809 ();
 FILLCELL_X4 FILLER_104_825 ();
 FILLCELL_X2 FILLER_104_829 ();
 FILLCELL_X1 FILLER_104_831 ();
 FILLCELL_X8 FILLER_104_839 ();
 FILLCELL_X4 FILLER_104_847 ();
 FILLCELL_X1 FILLER_104_851 ();
 FILLCELL_X4 FILLER_104_877 ();
 FILLCELL_X2 FILLER_104_903 ();
 FILLCELL_X8 FILLER_104_918 ();
 FILLCELL_X4 FILLER_104_926 ();
 FILLCELL_X2 FILLER_104_930 ();
 FILLCELL_X8 FILLER_104_941 ();
 FILLCELL_X4 FILLER_104_949 ();
 FILLCELL_X2 FILLER_104_953 ();
 FILLCELL_X1 FILLER_104_955 ();
 FILLCELL_X16 FILLER_104_972 ();
 FILLCELL_X4 FILLER_104_988 ();
 FILLCELL_X2 FILLER_104_992 ();
 FILLCELL_X1 FILLER_104_1010 ();
 FILLCELL_X2 FILLER_104_1018 ();
 FILLCELL_X1 FILLER_104_1023 ();
 FILLCELL_X2 FILLER_104_1042 ();
 FILLCELL_X1 FILLER_104_1044 ();
 FILLCELL_X8 FILLER_104_1066 ();
 FILLCELL_X4 FILLER_104_1074 ();
 FILLCELL_X1 FILLER_104_1088 ();
 FILLCELL_X2 FILLER_104_1110 ();
 FILLCELL_X8 FILLER_104_1123 ();
 FILLCELL_X4 FILLER_104_1131 ();
 FILLCELL_X2 FILLER_104_1145 ();
 FILLCELL_X1 FILLER_104_1172 ();
 FILLCELL_X8 FILLER_104_1180 ();
 FILLCELL_X2 FILLER_104_1188 ();
 FILLCELL_X1 FILLER_104_1190 ();
 FILLCELL_X8 FILLER_104_1194 ();
 FILLCELL_X4 FILLER_104_1202 ();
 FILLCELL_X2 FILLER_104_1206 ();
 FILLCELL_X1 FILLER_104_1208 ();
 FILLCELL_X16 FILLER_105_1 ();
 FILLCELL_X1 FILLER_105_17 ();
 FILLCELL_X32 FILLER_105_21 ();
 FILLCELL_X32 FILLER_105_53 ();
 FILLCELL_X16 FILLER_105_85 ();
 FILLCELL_X8 FILLER_105_101 ();
 FILLCELL_X1 FILLER_105_109 ();
 FILLCELL_X2 FILLER_105_123 ();
 FILLCELL_X1 FILLER_105_125 ();
 FILLCELL_X4 FILLER_105_161 ();
 FILLCELL_X2 FILLER_105_165 ();
 FILLCELL_X2 FILLER_105_174 ();
 FILLCELL_X1 FILLER_105_176 ();
 FILLCELL_X4 FILLER_105_187 ();
 FILLCELL_X2 FILLER_105_191 ();
 FILLCELL_X1 FILLER_105_193 ();
 FILLCELL_X4 FILLER_105_221 ();
 FILLCELL_X4 FILLER_105_238 ();
 FILLCELL_X2 FILLER_105_242 ();
 FILLCELL_X2 FILLER_105_256 ();
 FILLCELL_X32 FILLER_105_271 ();
 FILLCELL_X16 FILLER_105_303 ();
 FILLCELL_X4 FILLER_105_319 ();
 FILLCELL_X2 FILLER_105_323 ();
 FILLCELL_X1 FILLER_105_325 ();
 FILLCELL_X16 FILLER_105_336 ();
 FILLCELL_X2 FILLER_105_352 ();
 FILLCELL_X8 FILLER_105_363 ();
 FILLCELL_X4 FILLER_105_371 ();
 FILLCELL_X2 FILLER_105_375 ();
 FILLCELL_X8 FILLER_105_386 ();
 FILLCELL_X4 FILLER_105_394 ();
 FILLCELL_X2 FILLER_105_398 ();
 FILLCELL_X2 FILLER_105_422 ();
 FILLCELL_X2 FILLER_105_451 ();
 FILLCELL_X1 FILLER_105_453 ();
 FILLCELL_X16 FILLER_105_463 ();
 FILLCELL_X4 FILLER_105_479 ();
 FILLCELL_X2 FILLER_105_483 ();
 FILLCELL_X1 FILLER_105_485 ();
 FILLCELL_X1 FILLER_105_493 ();
 FILLCELL_X2 FILLER_105_523 ();
 FILLCELL_X2 FILLER_105_570 ();
 FILLCELL_X1 FILLER_105_572 ();
 FILLCELL_X2 FILLER_105_590 ();
 FILLCELL_X4 FILLER_105_595 ();
 FILLCELL_X1 FILLER_105_599 ();
 FILLCELL_X8 FILLER_105_611 ();
 FILLCELL_X8 FILLER_105_628 ();
 FILLCELL_X4 FILLER_105_636 ();
 FILLCELL_X1 FILLER_105_640 ();
 FILLCELL_X4 FILLER_105_653 ();
 FILLCELL_X1 FILLER_105_657 ();
 FILLCELL_X16 FILLER_105_665 ();
 FILLCELL_X2 FILLER_105_681 ();
 FILLCELL_X2 FILLER_105_690 ();
 FILLCELL_X1 FILLER_105_692 ();
 FILLCELL_X32 FILLER_105_697 ();
 FILLCELL_X8 FILLER_105_729 ();
 FILLCELL_X2 FILLER_105_737 ();
 FILLCELL_X4 FILLER_105_741 ();
 FILLCELL_X2 FILLER_105_745 ();
 FILLCELL_X1 FILLER_105_747 ();
 FILLCELL_X16 FILLER_105_768 ();
 FILLCELL_X8 FILLER_105_784 ();
 FILLCELL_X8 FILLER_105_798 ();
 FILLCELL_X2 FILLER_105_806 ();
 FILLCELL_X1 FILLER_105_808 ();
 FILLCELL_X8 FILLER_105_816 ();
 FILLCELL_X2 FILLER_105_824 ();
 FILLCELL_X4 FILLER_105_848 ();
 FILLCELL_X2 FILLER_105_852 ();
 FILLCELL_X2 FILLER_105_902 ();
 FILLCELL_X1 FILLER_105_904 ();
 FILLCELL_X1 FILLER_105_919 ();
 FILLCELL_X2 FILLER_105_929 ();
 FILLCELL_X1 FILLER_105_931 ();
 FILLCELL_X4 FILLER_105_949 ();
 FILLCELL_X2 FILLER_105_953 ();
 FILLCELL_X8 FILLER_105_979 ();
 FILLCELL_X2 FILLER_105_987 ();
 FILLCELL_X8 FILLER_105_1038 ();
 FILLCELL_X2 FILLER_105_1046 ();
 FILLCELL_X1 FILLER_105_1048 ();
 FILLCELL_X16 FILLER_105_1071 ();
 FILLCELL_X4 FILLER_105_1087 ();
 FILLCELL_X2 FILLER_105_1091 ();
 FILLCELL_X1 FILLER_105_1093 ();
 FILLCELL_X1 FILLER_105_1100 ();
 FILLCELL_X1 FILLER_105_1121 ();
 FILLCELL_X1 FILLER_105_1152 ();
 FILLCELL_X2 FILLER_105_1164 ();
 FILLCELL_X4 FILLER_105_1170 ();
 FILLCELL_X2 FILLER_105_1177 ();
 FILLCELL_X8 FILLER_105_1188 ();
 FILLCELL_X1 FILLER_105_1196 ();
 FILLCELL_X8 FILLER_105_1201 ();
 FILLCELL_X32 FILLER_106_1 ();
 FILLCELL_X32 FILLER_106_33 ();
 FILLCELL_X32 FILLER_106_65 ();
 FILLCELL_X8 FILLER_106_97 ();
 FILLCELL_X4 FILLER_106_105 ();
 FILLCELL_X4 FILLER_106_151 ();
 FILLCELL_X1 FILLER_106_155 ();
 FILLCELL_X4 FILLER_106_167 ();
 FILLCELL_X1 FILLER_106_171 ();
 FILLCELL_X2 FILLER_106_181 ();
 FILLCELL_X1 FILLER_106_192 ();
 FILLCELL_X2 FILLER_106_204 ();
 FILLCELL_X1 FILLER_106_210 ();
 FILLCELL_X1 FILLER_106_220 ();
 FILLCELL_X1 FILLER_106_226 ();
 FILLCELL_X1 FILLER_106_236 ();
 FILLCELL_X32 FILLER_106_268 ();
 FILLCELL_X16 FILLER_106_300 ();
 FILLCELL_X4 FILLER_106_316 ();
 FILLCELL_X2 FILLER_106_320 ();
 FILLCELL_X4 FILLER_106_329 ();
 FILLCELL_X2 FILLER_106_333 ();
 FILLCELL_X2 FILLER_106_352 ();
 FILLCELL_X1 FILLER_106_354 ();
 FILLCELL_X4 FILLER_106_358 ();
 FILLCELL_X2 FILLER_106_362 ();
 FILLCELL_X1 FILLER_106_364 ();
 FILLCELL_X4 FILLER_106_367 ();
 FILLCELL_X2 FILLER_106_371 ();
 FILLCELL_X4 FILLER_106_414 ();
 FILLCELL_X8 FILLER_106_425 ();
 FILLCELL_X4 FILLER_106_433 ();
 FILLCELL_X2 FILLER_106_437 ();
 FILLCELL_X8 FILLER_106_442 ();
 FILLCELL_X32 FILLER_106_467 ();
 FILLCELL_X4 FILLER_106_499 ();
 FILLCELL_X2 FILLER_106_503 ();
 FILLCELL_X2 FILLER_106_511 ();
 FILLCELL_X1 FILLER_106_533 ();
 FILLCELL_X2 FILLER_106_542 ();
 FILLCELL_X1 FILLER_106_544 ();
 FILLCELL_X8 FILLER_106_552 ();
 FILLCELL_X2 FILLER_106_560 ();
 FILLCELL_X1 FILLER_106_562 ();
 FILLCELL_X4 FILLER_106_585 ();
 FILLCELL_X1 FILLER_106_589 ();
 FILLCELL_X2 FILLER_106_608 ();
 FILLCELL_X1 FILLER_106_610 ();
 FILLCELL_X4 FILLER_106_627 ();
 FILLCELL_X8 FILLER_106_632 ();
 FILLCELL_X4 FILLER_106_640 ();
 FILLCELL_X2 FILLER_106_644 ();
 FILLCELL_X1 FILLER_106_650 ();
 FILLCELL_X2 FILLER_106_668 ();
 FILLCELL_X1 FILLER_106_670 ();
 FILLCELL_X2 FILLER_106_686 ();
 FILLCELL_X16 FILLER_106_709 ();
 FILLCELL_X8 FILLER_106_725 ();
 FILLCELL_X4 FILLER_106_750 ();
 FILLCELL_X16 FILLER_106_773 ();
 FILLCELL_X1 FILLER_106_789 ();
 FILLCELL_X4 FILLER_106_803 ();
 FILLCELL_X2 FILLER_106_807 ();
 FILLCELL_X2 FILLER_106_819 ();
 FILLCELL_X1 FILLER_106_821 ();
 FILLCELL_X2 FILLER_106_850 ();
 FILLCELL_X2 FILLER_106_860 ();
 FILLCELL_X1 FILLER_106_862 ();
 FILLCELL_X2 FILLER_106_870 ();
 FILLCELL_X2 FILLER_106_879 ();
 FILLCELL_X1 FILLER_106_906 ();
 FILLCELL_X1 FILLER_106_916 ();
 FILLCELL_X2 FILLER_106_924 ();
 FILLCELL_X2 FILLER_106_935 ();
 FILLCELL_X1 FILLER_106_937 ();
 FILLCELL_X2 FILLER_106_958 ();
 FILLCELL_X16 FILLER_106_977 ();
 FILLCELL_X8 FILLER_106_993 ();
 FILLCELL_X4 FILLER_106_1001 ();
 FILLCELL_X2 FILLER_106_1005 ();
 FILLCELL_X4 FILLER_106_1016 ();
 FILLCELL_X16 FILLER_106_1023 ();
 FILLCELL_X8 FILLER_106_1056 ();
 FILLCELL_X1 FILLER_106_1064 ();
 FILLCELL_X1 FILLER_106_1079 ();
 FILLCELL_X2 FILLER_106_1084 ();
 FILLCELL_X1 FILLER_106_1086 ();
 FILLCELL_X2 FILLER_106_1091 ();
 FILLCELL_X2 FILLER_106_1114 ();
 FILLCELL_X2 FILLER_106_1131 ();
 FILLCELL_X1 FILLER_106_1133 ();
 FILLCELL_X1 FILLER_106_1146 ();
 FILLCELL_X1 FILLER_106_1159 ();
 FILLCELL_X2 FILLER_106_1178 ();
 FILLCELL_X1 FILLER_106_1180 ();
 FILLCELL_X4 FILLER_106_1189 ();
 FILLCELL_X2 FILLER_106_1193 ();
 FILLCELL_X8 FILLER_106_1198 ();
 FILLCELL_X2 FILLER_106_1206 ();
 FILLCELL_X1 FILLER_106_1208 ();
 FILLCELL_X16 FILLER_107_1 ();
 FILLCELL_X8 FILLER_107_17 ();
 FILLCELL_X32 FILLER_107_28 ();
 FILLCELL_X32 FILLER_107_60 ();
 FILLCELL_X8 FILLER_107_92 ();
 FILLCELL_X1 FILLER_107_100 ();
 FILLCELL_X1 FILLER_107_114 ();
 FILLCELL_X2 FILLER_107_119 ();
 FILLCELL_X2 FILLER_107_148 ();
 FILLCELL_X1 FILLER_107_162 ();
 FILLCELL_X1 FILLER_107_169 ();
 FILLCELL_X2 FILLER_107_184 ();
 FILLCELL_X1 FILLER_107_206 ();
 FILLCELL_X1 FILLER_107_211 ();
 FILLCELL_X8 FILLER_107_215 ();
 FILLCELL_X1 FILLER_107_223 ();
 FILLCELL_X4 FILLER_107_235 ();
 FILLCELL_X2 FILLER_107_239 ();
 FILLCELL_X2 FILLER_107_250 ();
 FILLCELL_X2 FILLER_107_261 ();
 FILLCELL_X2 FILLER_107_269 ();
 FILLCELL_X2 FILLER_107_285 ();
 FILLCELL_X1 FILLER_107_287 ();
 FILLCELL_X4 FILLER_107_359 ();
 FILLCELL_X1 FILLER_107_363 ();
 FILLCELL_X4 FILLER_107_382 ();
 FILLCELL_X2 FILLER_107_386 ();
 FILLCELL_X8 FILLER_107_392 ();
 FILLCELL_X4 FILLER_107_400 ();
 FILLCELL_X1 FILLER_107_404 ();
 FILLCELL_X32 FILLER_107_421 ();
 FILLCELL_X32 FILLER_107_453 ();
 FILLCELL_X16 FILLER_107_485 ();
 FILLCELL_X4 FILLER_107_501 ();
 FILLCELL_X2 FILLER_107_505 ();
 FILLCELL_X1 FILLER_107_514 ();
 FILLCELL_X16 FILLER_107_529 ();
 FILLCELL_X8 FILLER_107_545 ();
 FILLCELL_X4 FILLER_107_553 ();
 FILLCELL_X1 FILLER_107_557 ();
 FILLCELL_X8 FILLER_107_561 ();
 FILLCELL_X2 FILLER_107_590 ();
 FILLCELL_X2 FILLER_107_604 ();
 FILLCELL_X1 FILLER_107_606 ();
 FILLCELL_X1 FILLER_107_614 ();
 FILLCELL_X2 FILLER_107_626 ();
 FILLCELL_X2 FILLER_107_635 ();
 FILLCELL_X2 FILLER_107_646 ();
 FILLCELL_X4 FILLER_107_661 ();
 FILLCELL_X2 FILLER_107_665 ();
 FILLCELL_X1 FILLER_107_667 ();
 FILLCELL_X4 FILLER_107_684 ();
 FILLCELL_X1 FILLER_107_688 ();
 FILLCELL_X2 FILLER_107_696 ();
 FILLCELL_X1 FILLER_107_698 ();
 FILLCELL_X32 FILLER_107_712 ();
 FILLCELL_X16 FILLER_107_744 ();
 FILLCELL_X8 FILLER_107_760 ();
 FILLCELL_X4 FILLER_107_768 ();
 FILLCELL_X1 FILLER_107_772 ();
 FILLCELL_X4 FILLER_107_780 ();
 FILLCELL_X1 FILLER_107_784 ();
 FILLCELL_X2 FILLER_107_814 ();
 FILLCELL_X1 FILLER_107_837 ();
 FILLCELL_X2 FILLER_107_842 ();
 FILLCELL_X2 FILLER_107_848 ();
 FILLCELL_X2 FILLER_107_855 ();
 FILLCELL_X4 FILLER_107_907 ();
 FILLCELL_X1 FILLER_107_911 ();
 FILLCELL_X1 FILLER_107_919 ();
 FILLCELL_X2 FILLER_107_927 ();
 FILLCELL_X8 FILLER_107_939 ();
 FILLCELL_X4 FILLER_107_947 ();
 FILLCELL_X8 FILLER_107_979 ();
 FILLCELL_X2 FILLER_107_987 ();
 FILLCELL_X2 FILLER_107_1000 ();
 FILLCELL_X1 FILLER_107_1002 ();
 FILLCELL_X2 FILLER_107_1017 ();
 FILLCELL_X1 FILLER_107_1019 ();
 FILLCELL_X2 FILLER_107_1040 ();
 FILLCELL_X1 FILLER_107_1042 ();
 FILLCELL_X1 FILLER_107_1093 ();
 FILLCELL_X2 FILLER_107_1154 ();
 FILLCELL_X2 FILLER_107_1166 ();
 FILLCELL_X16 FILLER_107_1181 ();
 FILLCELL_X8 FILLER_107_1197 ();
 FILLCELL_X4 FILLER_107_1205 ();
 FILLCELL_X32 FILLER_108_1 ();
 FILLCELL_X32 FILLER_108_33 ();
 FILLCELL_X32 FILLER_108_65 ();
 FILLCELL_X4 FILLER_108_97 ();
 FILLCELL_X2 FILLER_108_101 ();
 FILLCELL_X1 FILLER_108_134 ();
 FILLCELL_X4 FILLER_108_152 ();
 FILLCELL_X1 FILLER_108_156 ();
 FILLCELL_X4 FILLER_108_164 ();
 FILLCELL_X1 FILLER_108_168 ();
 FILLCELL_X2 FILLER_108_173 ();
 FILLCELL_X1 FILLER_108_180 ();
 FILLCELL_X4 FILLER_108_191 ();
 FILLCELL_X2 FILLER_108_195 ();
 FILLCELL_X1 FILLER_108_226 ();
 FILLCELL_X1 FILLER_108_240 ();
 FILLCELL_X1 FILLER_108_245 ();
 FILLCELL_X1 FILLER_108_254 ();
 FILLCELL_X16 FILLER_108_271 ();
 FILLCELL_X8 FILLER_108_287 ();
 FILLCELL_X1 FILLER_108_303 ();
 FILLCELL_X8 FILLER_108_317 ();
 FILLCELL_X4 FILLER_108_325 ();
 FILLCELL_X4 FILLER_108_336 ();
 FILLCELL_X1 FILLER_108_340 ();
 FILLCELL_X2 FILLER_108_345 ();
 FILLCELL_X4 FILLER_108_367 ();
 FILLCELL_X1 FILLER_108_371 ();
 FILLCELL_X8 FILLER_108_399 ();
 FILLCELL_X4 FILLER_108_407 ();
 FILLCELL_X1 FILLER_108_411 ();
 FILLCELL_X1 FILLER_108_416 ();
 FILLCELL_X1 FILLER_108_423 ();
 FILLCELL_X32 FILLER_108_444 ();
 FILLCELL_X32 FILLER_108_476 ();
 FILLCELL_X2 FILLER_108_508 ();
 FILLCELL_X1 FILLER_108_510 ();
 FILLCELL_X2 FILLER_108_521 ();
 FILLCELL_X1 FILLER_108_523 ();
 FILLCELL_X8 FILLER_108_534 ();
 FILLCELL_X4 FILLER_108_546 ();
 FILLCELL_X1 FILLER_108_550 ();
 FILLCELL_X8 FILLER_108_571 ();
 FILLCELL_X2 FILLER_108_589 ();
 FILLCELL_X4 FILLER_108_595 ();
 FILLCELL_X2 FILLER_108_599 ();
 FILLCELL_X4 FILLER_108_611 ();
 FILLCELL_X2 FILLER_108_615 ();
 FILLCELL_X1 FILLER_108_617 ();
 FILLCELL_X8 FILLER_108_622 ();
 FILLCELL_X1 FILLER_108_630 ();
 FILLCELL_X2 FILLER_108_636 ();
 FILLCELL_X1 FILLER_108_638 ();
 FILLCELL_X1 FILLER_108_651 ();
 FILLCELL_X1 FILLER_108_662 ();
 FILLCELL_X4 FILLER_108_691 ();
 FILLCELL_X2 FILLER_108_695 ();
 FILLCELL_X1 FILLER_108_697 ();
 FILLCELL_X32 FILLER_108_711 ();
 FILLCELL_X32 FILLER_108_743 ();
 FILLCELL_X8 FILLER_108_775 ();
 FILLCELL_X2 FILLER_108_794 ();
 FILLCELL_X4 FILLER_108_804 ();
 FILLCELL_X2 FILLER_108_812 ();
 FILLCELL_X1 FILLER_108_814 ();
 FILLCELL_X4 FILLER_108_819 ();
 FILLCELL_X1 FILLER_108_823 ();
 FILLCELL_X8 FILLER_108_828 ();
 FILLCELL_X4 FILLER_108_836 ();
 FILLCELL_X2 FILLER_108_840 ();
 FILLCELL_X1 FILLER_108_842 ();
 FILLCELL_X8 FILLER_108_850 ();
 FILLCELL_X2 FILLER_108_861 ();
 FILLCELL_X1 FILLER_108_872 ();
 FILLCELL_X1 FILLER_108_909 ();
 FILLCELL_X2 FILLER_108_919 ();
 FILLCELL_X1 FILLER_108_921 ();
 FILLCELL_X8 FILLER_108_945 ();
 FILLCELL_X4 FILLER_108_953 ();
 FILLCELL_X32 FILLER_108_960 ();
 FILLCELL_X8 FILLER_108_992 ();
 FILLCELL_X4 FILLER_108_1000 ();
 FILLCELL_X2 FILLER_108_1004 ();
 FILLCELL_X1 FILLER_108_1006 ();
 FILLCELL_X4 FILLER_108_1020 ();
 FILLCELL_X2 FILLER_108_1024 ();
 FILLCELL_X1 FILLER_108_1026 ();
 FILLCELL_X2 FILLER_108_1060 ();
 FILLCELL_X1 FILLER_108_1062 ();
 FILLCELL_X2 FILLER_108_1080 ();
 FILLCELL_X1 FILLER_108_1082 ();
 FILLCELL_X16 FILLER_108_1090 ();
 FILLCELL_X2 FILLER_108_1106 ();
 FILLCELL_X2 FILLER_108_1111 ();
 FILLCELL_X8 FILLER_108_1142 ();
 FILLCELL_X1 FILLER_108_1167 ();
 FILLCELL_X1 FILLER_108_1172 ();
 FILLCELL_X2 FILLER_108_1177 ();
 FILLCELL_X8 FILLER_108_1185 ();
 FILLCELL_X1 FILLER_108_1193 ();
 FILLCELL_X8 FILLER_108_1197 ();
 FILLCELL_X4 FILLER_108_1205 ();
 FILLCELL_X2 FILLER_109_1 ();
 FILLCELL_X32 FILLER_109_6 ();
 FILLCELL_X32 FILLER_109_38 ();
 FILLCELL_X32 FILLER_109_70 ();
 FILLCELL_X4 FILLER_109_102 ();
 FILLCELL_X1 FILLER_109_110 ();
 FILLCELL_X1 FILLER_109_127 ();
 FILLCELL_X1 FILLER_109_143 ();
 FILLCELL_X1 FILLER_109_149 ();
 FILLCELL_X1 FILLER_109_155 ();
 FILLCELL_X8 FILLER_109_172 ();
 FILLCELL_X4 FILLER_109_180 ();
 FILLCELL_X8 FILLER_109_195 ();
 FILLCELL_X2 FILLER_109_203 ();
 FILLCELL_X1 FILLER_109_205 ();
 FILLCELL_X1 FILLER_109_241 ();
 FILLCELL_X1 FILLER_109_254 ();
 FILLCELL_X32 FILLER_109_273 ();
 FILLCELL_X2 FILLER_109_305 ();
 FILLCELL_X2 FILLER_109_328 ();
 FILLCELL_X8 FILLER_109_335 ();
 FILLCELL_X1 FILLER_109_343 ();
 FILLCELL_X1 FILLER_109_349 ();
 FILLCELL_X4 FILLER_109_357 ();
 FILLCELL_X2 FILLER_109_375 ();
 FILLCELL_X4 FILLER_109_383 ();
 FILLCELL_X1 FILLER_109_387 ();
 FILLCELL_X8 FILLER_109_392 ();
 FILLCELL_X4 FILLER_109_400 ();
 FILLCELL_X2 FILLER_109_408 ();
 FILLCELL_X1 FILLER_109_410 ();
 FILLCELL_X1 FILLER_109_422 ();
 FILLCELL_X8 FILLER_109_434 ();
 FILLCELL_X1 FILLER_109_442 ();
 FILLCELL_X32 FILLER_109_457 ();
 FILLCELL_X16 FILLER_109_489 ();
 FILLCELL_X2 FILLER_109_505 ();
 FILLCELL_X8 FILLER_109_517 ();
 FILLCELL_X2 FILLER_109_531 ();
 FILLCELL_X1 FILLER_109_536 ();
 FILLCELL_X1 FILLER_109_542 ();
 FILLCELL_X16 FILLER_109_555 ();
 FILLCELL_X8 FILLER_109_571 ();
 FILLCELL_X16 FILLER_109_590 ();
 FILLCELL_X1 FILLER_109_606 ();
 FILLCELL_X1 FILLER_109_611 ();
 FILLCELL_X8 FILLER_109_616 ();
 FILLCELL_X4 FILLER_109_624 ();
 FILLCELL_X1 FILLER_109_628 ();
 FILLCELL_X8 FILLER_109_633 ();
 FILLCELL_X8 FILLER_109_652 ();
 FILLCELL_X1 FILLER_109_670 ();
 FILLCELL_X2 FILLER_109_676 ();
 FILLCELL_X4 FILLER_109_691 ();
 FILLCELL_X1 FILLER_109_695 ();
 FILLCELL_X2 FILLER_109_703 ();
 FILLCELL_X32 FILLER_109_718 ();
 FILLCELL_X8 FILLER_109_750 ();
 FILLCELL_X4 FILLER_109_758 ();
 FILLCELL_X1 FILLER_109_791 ();
 FILLCELL_X4 FILLER_109_801 ();
 FILLCELL_X2 FILLER_109_805 ();
 FILLCELL_X1 FILLER_109_807 ();
 FILLCELL_X8 FILLER_109_812 ();
 FILLCELL_X2 FILLER_109_820 ();
 FILLCELL_X1 FILLER_109_822 ();
 FILLCELL_X4 FILLER_109_831 ();
 FILLCELL_X1 FILLER_109_864 ();
 FILLCELL_X2 FILLER_109_875 ();
 FILLCELL_X1 FILLER_109_903 ();
 FILLCELL_X1 FILLER_109_915 ();
 FILLCELL_X16 FILLER_109_936 ();
 FILLCELL_X8 FILLER_109_952 ();
 FILLCELL_X4 FILLER_109_960 ();
 FILLCELL_X2 FILLER_109_964 ();
 FILLCELL_X8 FILLER_109_983 ();
 FILLCELL_X4 FILLER_109_991 ();
 FILLCELL_X2 FILLER_109_995 ();
 FILLCELL_X4 FILLER_109_1004 ();
 FILLCELL_X2 FILLER_109_1019 ();
 FILLCELL_X1 FILLER_109_1021 ();
 FILLCELL_X1 FILLER_109_1037 ();
 FILLCELL_X1 FILLER_109_1061 ();
 FILLCELL_X2 FILLER_109_1072 ();
 FILLCELL_X1 FILLER_109_1074 ();
 FILLCELL_X1 FILLER_109_1104 ();
 FILLCELL_X4 FILLER_109_1112 ();
 FILLCELL_X2 FILLER_109_1116 ();
 FILLCELL_X1 FILLER_109_1118 ();
 FILLCELL_X8 FILLER_109_1124 ();
 FILLCELL_X2 FILLER_109_1132 ();
 FILLCELL_X1 FILLER_109_1134 ();
 FILLCELL_X4 FILLER_109_1141 ();
 FILLCELL_X1 FILLER_109_1145 ();
 FILLCELL_X2 FILLER_109_1150 ();
 FILLCELL_X1 FILLER_109_1158 ();
 FILLCELL_X2 FILLER_109_1164 ();
 FILLCELL_X1 FILLER_109_1166 ();
 FILLCELL_X16 FILLER_109_1185 ();
 FILLCELL_X8 FILLER_109_1201 ();
 FILLCELL_X32 FILLER_110_1 ();
 FILLCELL_X32 FILLER_110_33 ();
 FILLCELL_X32 FILLER_110_65 ();
 FILLCELL_X8 FILLER_110_97 ();
 FILLCELL_X4 FILLER_110_125 ();
 FILLCELL_X2 FILLER_110_133 ();
 FILLCELL_X1 FILLER_110_135 ();
 FILLCELL_X1 FILLER_110_143 ();
 FILLCELL_X2 FILLER_110_151 ();
 FILLCELL_X4 FILLER_110_155 ();
 FILLCELL_X2 FILLER_110_159 ();
 FILLCELL_X2 FILLER_110_172 ();
 FILLCELL_X2 FILLER_110_200 ();
 FILLCELL_X1 FILLER_110_202 ();
 FILLCELL_X2 FILLER_110_210 ();
 FILLCELL_X8 FILLER_110_232 ();
 FILLCELL_X2 FILLER_110_240 ();
 FILLCELL_X1 FILLER_110_266 ();
 FILLCELL_X32 FILLER_110_270 ();
 FILLCELL_X2 FILLER_110_302 ();
 FILLCELL_X2 FILLER_110_318 ();
 FILLCELL_X1 FILLER_110_320 ();
 FILLCELL_X1 FILLER_110_358 ();
 FILLCELL_X2 FILLER_110_384 ();
 FILLCELL_X2 FILLER_110_412 ();
 FILLCELL_X4 FILLER_110_418 ();
 FILLCELL_X4 FILLER_110_440 ();
 FILLCELL_X32 FILLER_110_451 ();
 FILLCELL_X8 FILLER_110_483 ();
 FILLCELL_X2 FILLER_110_491 ();
 FILLCELL_X2 FILLER_110_500 ();
 FILLCELL_X1 FILLER_110_513 ();
 FILLCELL_X1 FILLER_110_537 ();
 FILLCELL_X1 FILLER_110_545 ();
 FILLCELL_X1 FILLER_110_550 ();
 FILLCELL_X1 FILLER_110_556 ();
 FILLCELL_X4 FILLER_110_563 ();
 FILLCELL_X1 FILLER_110_567 ();
 FILLCELL_X8 FILLER_110_572 ();
 FILLCELL_X4 FILLER_110_580 ();
 FILLCELL_X2 FILLER_110_584 ();
 FILLCELL_X1 FILLER_110_586 ();
 FILLCELL_X2 FILLER_110_590 ();
 FILLCELL_X1 FILLER_110_651 ();
 FILLCELL_X2 FILLER_110_672 ();
 FILLCELL_X1 FILLER_110_696 ();
 FILLCELL_X8 FILLER_110_706 ();
 FILLCELL_X32 FILLER_110_723 ();
 FILLCELL_X8 FILLER_110_755 ();
 FILLCELL_X1 FILLER_110_763 ();
 FILLCELL_X1 FILLER_110_768 ();
 FILLCELL_X2 FILLER_110_772 ();
 FILLCELL_X1 FILLER_110_774 ();
 FILLCELL_X2 FILLER_110_779 ();
 FILLCELL_X1 FILLER_110_781 ();
 FILLCELL_X4 FILLER_110_800 ();
 FILLCELL_X2 FILLER_110_814 ();
 FILLCELL_X2 FILLER_110_827 ();
 FILLCELL_X2 FILLER_110_833 ();
 FILLCELL_X2 FILLER_110_842 ();
 FILLCELL_X8 FILLER_110_882 ();
 FILLCELL_X2 FILLER_110_890 ();
 FILLCELL_X1 FILLER_110_892 ();
 FILLCELL_X4 FILLER_110_921 ();
 FILLCELL_X2 FILLER_110_937 ();
 FILLCELL_X2 FILLER_110_973 ();
 FILLCELL_X16 FILLER_110_982 ();
 FILLCELL_X1 FILLER_110_998 ();
 FILLCELL_X1 FILLER_110_1008 ();
 FILLCELL_X4 FILLER_110_1016 ();
 FILLCELL_X2 FILLER_110_1020 ();
 FILLCELL_X1 FILLER_110_1040 ();
 FILLCELL_X8 FILLER_110_1079 ();
 FILLCELL_X1 FILLER_110_1087 ();
 FILLCELL_X4 FILLER_110_1092 ();
 FILLCELL_X2 FILLER_110_1096 ();
 FILLCELL_X1 FILLER_110_1098 ();
 FILLCELL_X4 FILLER_110_1113 ();
 FILLCELL_X1 FILLER_110_1117 ();
 FILLCELL_X2 FILLER_110_1121 ();
 FILLCELL_X2 FILLER_110_1131 ();
 FILLCELL_X4 FILLER_110_1141 ();
 FILLCELL_X2 FILLER_110_1145 ();
 FILLCELL_X1 FILLER_110_1147 ();
 FILLCELL_X2 FILLER_110_1178 ();
 FILLCELL_X1 FILLER_110_1190 ();
 FILLCELL_X8 FILLER_110_1198 ();
 FILLCELL_X2 FILLER_110_1206 ();
 FILLCELL_X1 FILLER_110_1208 ();
 FILLCELL_X8 FILLER_111_1 ();
 FILLCELL_X4 FILLER_111_9 ();
 FILLCELL_X2 FILLER_111_13 ();
 FILLCELL_X32 FILLER_111_19 ();
 FILLCELL_X32 FILLER_111_51 ();
 FILLCELL_X16 FILLER_111_83 ();
 FILLCELL_X4 FILLER_111_99 ();
 FILLCELL_X2 FILLER_111_117 ();
 FILLCELL_X1 FILLER_111_133 ();
 FILLCELL_X4 FILLER_111_156 ();
 FILLCELL_X1 FILLER_111_168 ();
 FILLCELL_X8 FILLER_111_177 ();
 FILLCELL_X4 FILLER_111_185 ();
 FILLCELL_X1 FILLER_111_189 ();
 FILLCELL_X4 FILLER_111_201 ();
 FILLCELL_X2 FILLER_111_205 ();
 FILLCELL_X1 FILLER_111_207 ();
 FILLCELL_X4 FILLER_111_215 ();
 FILLCELL_X1 FILLER_111_219 ();
 FILLCELL_X1 FILLER_111_238 ();
 FILLCELL_X1 FILLER_111_243 ();
 FILLCELL_X1 FILLER_111_252 ();
 FILLCELL_X8 FILLER_111_258 ();
 FILLCELL_X2 FILLER_111_266 ();
 FILLCELL_X32 FILLER_111_272 ();
 FILLCELL_X4 FILLER_111_304 ();
 FILLCELL_X2 FILLER_111_308 ();
 FILLCELL_X4 FILLER_111_326 ();
 FILLCELL_X2 FILLER_111_330 ();
 FILLCELL_X1 FILLER_111_341 ();
 FILLCELL_X1 FILLER_111_361 ();
 FILLCELL_X2 FILLER_111_397 ();
 FILLCELL_X1 FILLER_111_399 ();
 FILLCELL_X2 FILLER_111_405 ();
 FILLCELL_X1 FILLER_111_407 ();
 FILLCELL_X2 FILLER_111_424 ();
 FILLCELL_X1 FILLER_111_426 ();
 FILLCELL_X4 FILLER_111_432 ();
 FILLCELL_X2 FILLER_111_436 ();
 FILLCELL_X4 FILLER_111_445 ();
 FILLCELL_X32 FILLER_111_465 ();
 FILLCELL_X2 FILLER_111_497 ();
 FILLCELL_X2 FILLER_111_510 ();
 FILLCELL_X8 FILLER_111_516 ();
 FILLCELL_X2 FILLER_111_524 ();
 FILLCELL_X1 FILLER_111_530 ();
 FILLCELL_X8 FILLER_111_534 ();
 FILLCELL_X1 FILLER_111_542 ();
 FILLCELL_X8 FILLER_111_554 ();
 FILLCELL_X4 FILLER_111_562 ();
 FILLCELL_X2 FILLER_111_566 ();
 FILLCELL_X1 FILLER_111_568 ();
 FILLCELL_X1 FILLER_111_580 ();
 FILLCELL_X1 FILLER_111_584 ();
 FILLCELL_X2 FILLER_111_596 ();
 FILLCELL_X1 FILLER_111_603 ();
 FILLCELL_X2 FILLER_111_622 ();
 FILLCELL_X4 FILLER_111_636 ();
 FILLCELL_X2 FILLER_111_640 ();
 FILLCELL_X1 FILLER_111_642 ();
 FILLCELL_X4 FILLER_111_647 ();
 FILLCELL_X1 FILLER_111_651 ();
 FILLCELL_X16 FILLER_111_659 ();
 FILLCELL_X8 FILLER_111_675 ();
 FILLCELL_X1 FILLER_111_683 ();
 FILLCELL_X2 FILLER_111_691 ();
 FILLCELL_X1 FILLER_111_693 ();
 FILLCELL_X32 FILLER_111_739 ();
 FILLCELL_X4 FILLER_111_828 ();
 FILLCELL_X1 FILLER_111_832 ();
 FILLCELL_X2 FILLER_111_838 ();
 FILLCELL_X2 FILLER_111_863 ();
 FILLCELL_X1 FILLER_111_865 ();
 FILLCELL_X1 FILLER_111_880 ();
 FILLCELL_X2 FILLER_111_884 ();
 FILLCELL_X1 FILLER_111_886 ();
 FILLCELL_X2 FILLER_111_935 ();
 FILLCELL_X8 FILLER_111_944 ();
 FILLCELL_X4 FILLER_111_952 ();
 FILLCELL_X2 FILLER_111_956 ();
 FILLCELL_X4 FILLER_111_983 ();
 FILLCELL_X2 FILLER_111_987 ();
 FILLCELL_X1 FILLER_111_989 ();
 FILLCELL_X2 FILLER_111_1006 ();
 FILLCELL_X2 FILLER_111_1021 ();
 FILLCELL_X2 FILLER_111_1054 ();
 FILLCELL_X2 FILLER_111_1093 ();
 FILLCELL_X1 FILLER_111_1095 ();
 FILLCELL_X2 FILLER_111_1099 ();
 FILLCELL_X8 FILLER_111_1107 ();
 FILLCELL_X2 FILLER_111_1115 ();
 FILLCELL_X4 FILLER_111_1123 ();
 FILLCELL_X2 FILLER_111_1127 ();
 FILLCELL_X1 FILLER_111_1129 ();
 FILLCELL_X16 FILLER_111_1139 ();
 FILLCELL_X4 FILLER_111_1159 ();
 FILLCELL_X1 FILLER_111_1163 ();
 FILLCELL_X8 FILLER_111_1198 ();
 FILLCELL_X2 FILLER_111_1206 ();
 FILLCELL_X1 FILLER_111_1208 ();
 FILLCELL_X32 FILLER_112_1 ();
 FILLCELL_X32 FILLER_112_33 ();
 FILLCELL_X32 FILLER_112_65 ();
 FILLCELL_X8 FILLER_112_97 ();
 FILLCELL_X4 FILLER_112_105 ();
 FILLCELL_X1 FILLER_112_120 ();
 FILLCELL_X16 FILLER_112_147 ();
 FILLCELL_X1 FILLER_112_163 ();
 FILLCELL_X1 FILLER_112_171 ();
 FILLCELL_X1 FILLER_112_181 ();
 FILLCELL_X8 FILLER_112_187 ();
 FILLCELL_X1 FILLER_112_195 ();
 FILLCELL_X2 FILLER_112_199 ();
 FILLCELL_X1 FILLER_112_201 ();
 FILLCELL_X4 FILLER_112_210 ();
 FILLCELL_X2 FILLER_112_214 ();
 FILLCELL_X2 FILLER_112_227 ();
 FILLCELL_X1 FILLER_112_229 ();
 FILLCELL_X16 FILLER_112_273 ();
 FILLCELL_X8 FILLER_112_289 ();
 FILLCELL_X1 FILLER_112_297 ();
 FILLCELL_X1 FILLER_112_330 ();
 FILLCELL_X4 FILLER_112_342 ();
 FILLCELL_X2 FILLER_112_346 ();
 FILLCELL_X2 FILLER_112_356 ();
 FILLCELL_X1 FILLER_112_367 ();
 FILLCELL_X2 FILLER_112_378 ();
 FILLCELL_X1 FILLER_112_394 ();
 FILLCELL_X1 FILLER_112_419 ();
 FILLCELL_X2 FILLER_112_428 ();
 FILLCELL_X32 FILLER_112_450 ();
 FILLCELL_X8 FILLER_112_482 ();
 FILLCELL_X4 FILLER_112_490 ();
 FILLCELL_X2 FILLER_112_494 ();
 FILLCELL_X1 FILLER_112_496 ();
 FILLCELL_X8 FILLER_112_521 ();
 FILLCELL_X2 FILLER_112_529 ();
 FILLCELL_X1 FILLER_112_531 ();
 FILLCELL_X8 FILLER_112_552 ();
 FILLCELL_X1 FILLER_112_560 ();
 FILLCELL_X1 FILLER_112_568 ();
 FILLCELL_X4 FILLER_112_576 ();
 FILLCELL_X1 FILLER_112_580 ();
 FILLCELL_X1 FILLER_112_590 ();
 FILLCELL_X16 FILLER_112_615 ();
 FILLCELL_X4 FILLER_112_645 ();
 FILLCELL_X2 FILLER_112_649 ();
 FILLCELL_X1 FILLER_112_658 ();
 FILLCELL_X1 FILLER_112_688 ();
 FILLCELL_X4 FILLER_112_702 ();
 FILLCELL_X2 FILLER_112_706 ();
 FILLCELL_X32 FILLER_112_721 ();
 FILLCELL_X1 FILLER_112_753 ();
 FILLCELL_X2 FILLER_112_767 ();
 FILLCELL_X8 FILLER_112_794 ();
 FILLCELL_X4 FILLER_112_802 ();
 FILLCELL_X4 FILLER_112_810 ();
 FILLCELL_X2 FILLER_112_830 ();
 FILLCELL_X1 FILLER_112_832 ();
 FILLCELL_X4 FILLER_112_845 ();
 FILLCELL_X4 FILLER_112_852 ();
 FILLCELL_X2 FILLER_112_856 ();
 FILLCELL_X2 FILLER_112_869 ();
 FILLCELL_X1 FILLER_112_886 ();
 FILLCELL_X8 FILLER_112_895 ();
 FILLCELL_X2 FILLER_112_903 ();
 FILLCELL_X1 FILLER_112_905 ();
 FILLCELL_X32 FILLER_112_947 ();
 FILLCELL_X16 FILLER_112_979 ();
 FILLCELL_X8 FILLER_112_995 ();
 FILLCELL_X4 FILLER_112_1010 ();
 FILLCELL_X2 FILLER_112_1014 ();
 FILLCELL_X1 FILLER_112_1041 ();
 FILLCELL_X2 FILLER_112_1053 ();
 FILLCELL_X1 FILLER_112_1073 ();
 FILLCELL_X2 FILLER_112_1079 ();
 FILLCELL_X16 FILLER_112_1084 ();
 FILLCELL_X8 FILLER_112_1104 ();
 FILLCELL_X2 FILLER_112_1112 ();
 FILLCELL_X1 FILLER_112_1114 ();
 FILLCELL_X8 FILLER_112_1123 ();
 FILLCELL_X1 FILLER_112_1131 ();
 FILLCELL_X1 FILLER_112_1139 ();
 FILLCELL_X16 FILLER_112_1154 ();
 FILLCELL_X4 FILLER_112_1170 ();
 FILLCELL_X2 FILLER_112_1174 ();
 FILLCELL_X1 FILLER_112_1176 ();
 FILLCELL_X4 FILLER_112_1202 ();
 FILLCELL_X2 FILLER_112_1206 ();
 FILLCELL_X1 FILLER_112_1208 ();
 FILLCELL_X32 FILLER_113_1 ();
 FILLCELL_X32 FILLER_113_33 ();
 FILLCELL_X32 FILLER_113_65 ();
 FILLCELL_X8 FILLER_113_97 ();
 FILLCELL_X2 FILLER_113_105 ();
 FILLCELL_X1 FILLER_113_107 ();
 FILLCELL_X4 FILLER_113_112 ();
 FILLCELL_X1 FILLER_113_116 ();
 FILLCELL_X1 FILLER_113_130 ();
 FILLCELL_X1 FILLER_113_134 ();
 FILLCELL_X4 FILLER_113_149 ();
 FILLCELL_X2 FILLER_113_153 ();
 FILLCELL_X8 FILLER_113_168 ();
 FILLCELL_X2 FILLER_113_180 ();
 FILLCELL_X2 FILLER_113_186 ();
 FILLCELL_X2 FILLER_113_219 ();
 FILLCELL_X1 FILLER_113_221 ();
 FILLCELL_X2 FILLER_113_227 ();
 FILLCELL_X1 FILLER_113_234 ();
 FILLCELL_X2 FILLER_113_238 ();
 FILLCELL_X1 FILLER_113_240 ();
 FILLCELL_X2 FILLER_113_245 ();
 FILLCELL_X1 FILLER_113_247 ();
 FILLCELL_X1 FILLER_113_252 ();
 FILLCELL_X2 FILLER_113_256 ();
 FILLCELL_X1 FILLER_113_258 ();
 FILLCELL_X2 FILLER_113_262 ();
 FILLCELL_X16 FILLER_113_271 ();
 FILLCELL_X8 FILLER_113_287 ();
 FILLCELL_X2 FILLER_113_356 ();
 FILLCELL_X1 FILLER_113_358 ();
 FILLCELL_X2 FILLER_113_385 ();
 FILLCELL_X4 FILLER_113_394 ();
 FILLCELL_X1 FILLER_113_398 ();
 FILLCELL_X2 FILLER_113_419 ();
 FILLCELL_X4 FILLER_113_425 ();
 FILLCELL_X1 FILLER_113_429 ();
 FILLCELL_X1 FILLER_113_434 ();
 FILLCELL_X32 FILLER_113_457 ();
 FILLCELL_X8 FILLER_113_489 ();
 FILLCELL_X4 FILLER_113_497 ();
 FILLCELL_X1 FILLER_113_501 ();
 FILLCELL_X1 FILLER_113_511 ();
 FILLCELL_X8 FILLER_113_528 ();
 FILLCELL_X2 FILLER_113_536 ();
 FILLCELL_X1 FILLER_113_538 ();
 FILLCELL_X1 FILLER_113_550 ();
 FILLCELL_X1 FILLER_113_557 ();
 FILLCELL_X2 FILLER_113_562 ();
 FILLCELL_X1 FILLER_113_571 ();
 FILLCELL_X1 FILLER_113_576 ();
 FILLCELL_X2 FILLER_113_582 ();
 FILLCELL_X1 FILLER_113_584 ();
 FILLCELL_X16 FILLER_113_592 ();
 FILLCELL_X4 FILLER_113_615 ();
 FILLCELL_X2 FILLER_113_619 ();
 FILLCELL_X2 FILLER_113_635 ();
 FILLCELL_X1 FILLER_113_637 ();
 FILLCELL_X8 FILLER_113_678 ();
 FILLCELL_X2 FILLER_113_686 ();
 FILLCELL_X2 FILLER_113_705 ();
 FILLCELL_X1 FILLER_113_707 ();
 FILLCELL_X16 FILLER_113_728 ();
 FILLCELL_X8 FILLER_113_744 ();
 FILLCELL_X2 FILLER_113_752 ();
 FILLCELL_X1 FILLER_113_754 ();
 FILLCELL_X2 FILLER_113_773 ();
 FILLCELL_X2 FILLER_113_784 ();
 FILLCELL_X1 FILLER_113_786 ();
 FILLCELL_X1 FILLER_113_798 ();
 FILLCELL_X2 FILLER_113_810 ();
 FILLCELL_X1 FILLER_113_812 ();
 FILLCELL_X4 FILLER_113_821 ();
 FILLCELL_X8 FILLER_113_839 ();
 FILLCELL_X1 FILLER_113_847 ();
 FILLCELL_X4 FILLER_113_853 ();
 FILLCELL_X1 FILLER_113_857 ();
 FILLCELL_X1 FILLER_113_862 ();
 FILLCELL_X1 FILLER_113_867 ();
 FILLCELL_X4 FILLER_113_877 ();
 FILLCELL_X2 FILLER_113_881 ();
 FILLCELL_X1 FILLER_113_883 ();
 FILLCELL_X2 FILLER_113_888 ();
 FILLCELL_X2 FILLER_113_893 ();
 FILLCELL_X1 FILLER_113_895 ();
 FILLCELL_X2 FILLER_113_925 ();
 FILLCELL_X2 FILLER_113_930 ();
 FILLCELL_X16 FILLER_113_949 ();
 FILLCELL_X8 FILLER_113_965 ();
 FILLCELL_X1 FILLER_113_997 ();
 FILLCELL_X2 FILLER_113_1005 ();
 FILLCELL_X4 FILLER_113_1014 ();
 FILLCELL_X1 FILLER_113_1036 ();
 FILLCELL_X2 FILLER_113_1048 ();
 FILLCELL_X1 FILLER_113_1091 ();
 FILLCELL_X1 FILLER_113_1106 ();
 FILLCELL_X4 FILLER_113_1117 ();
 FILLCELL_X2 FILLER_113_1121 ();
 FILLCELL_X8 FILLER_113_1140 ();
 FILLCELL_X2 FILLER_113_1148 ();
 FILLCELL_X8 FILLER_113_1154 ();
 FILLCELL_X2 FILLER_113_1162 ();
 FILLCELL_X1 FILLER_113_1164 ();
 FILLCELL_X1 FILLER_113_1178 ();
 FILLCELL_X4 FILLER_113_1183 ();
 FILLCELL_X2 FILLER_113_1187 ();
 FILLCELL_X1 FILLER_113_1189 ();
 FILLCELL_X16 FILLER_113_1193 ();
 FILLCELL_X8 FILLER_114_1 ();
 FILLCELL_X4 FILLER_114_9 ();
 FILLCELL_X32 FILLER_114_16 ();
 FILLCELL_X32 FILLER_114_48 ();
 FILLCELL_X16 FILLER_114_80 ();
 FILLCELL_X8 FILLER_114_96 ();
 FILLCELL_X2 FILLER_114_104 ();
 FILLCELL_X1 FILLER_114_106 ();
 FILLCELL_X4 FILLER_114_116 ();
 FILLCELL_X2 FILLER_114_120 ();
 FILLCELL_X1 FILLER_114_126 ();
 FILLCELL_X1 FILLER_114_142 ();
 FILLCELL_X1 FILLER_114_150 ();
 FILLCELL_X1 FILLER_114_156 ();
 FILLCELL_X4 FILLER_114_168 ();
 FILLCELL_X1 FILLER_114_172 ();
 FILLCELL_X2 FILLER_114_178 ();
 FILLCELL_X2 FILLER_114_241 ();
 FILLCELL_X1 FILLER_114_243 ();
 FILLCELL_X4 FILLER_114_253 ();
 FILLCELL_X8 FILLER_114_267 ();
 FILLCELL_X2 FILLER_114_275 ();
 FILLCELL_X1 FILLER_114_277 ();
 FILLCELL_X2 FILLER_114_302 ();
 FILLCELL_X2 FILLER_114_334 ();
 FILLCELL_X2 FILLER_114_350 ();
 FILLCELL_X1 FILLER_114_352 ();
 FILLCELL_X1 FILLER_114_360 ();
 FILLCELL_X4 FILLER_114_367 ();
 FILLCELL_X1 FILLER_114_402 ();
 FILLCELL_X4 FILLER_114_407 ();
 FILLCELL_X2 FILLER_114_411 ();
 FILLCELL_X1 FILLER_114_413 ();
 FILLCELL_X4 FILLER_114_418 ();
 FILLCELL_X2 FILLER_114_433 ();
 FILLCELL_X1 FILLER_114_448 ();
 FILLCELL_X32 FILLER_114_456 ();
 FILLCELL_X16 FILLER_114_488 ();
 FILLCELL_X4 FILLER_114_504 ();
 FILLCELL_X4 FILLER_114_513 ();
 FILLCELL_X2 FILLER_114_517 ();
 FILLCELL_X4 FILLER_114_524 ();
 FILLCELL_X2 FILLER_114_538 ();
 FILLCELL_X2 FILLER_114_544 ();
 FILLCELL_X1 FILLER_114_546 ();
 FILLCELL_X4 FILLER_114_558 ();
 FILLCELL_X2 FILLER_114_562 ();
 FILLCELL_X8 FILLER_114_583 ();
 FILLCELL_X8 FILLER_114_598 ();
 FILLCELL_X2 FILLER_114_606 ();
 FILLCELL_X1 FILLER_114_608 ();
 FILLCELL_X1 FILLER_114_616 ();
 FILLCELL_X4 FILLER_114_627 ();
 FILLCELL_X4 FILLER_114_632 ();
 FILLCELL_X1 FILLER_114_636 ();
 FILLCELL_X2 FILLER_114_644 ();
 FILLCELL_X2 FILLER_114_649 ();
 FILLCELL_X8 FILLER_114_676 ();
 FILLCELL_X4 FILLER_114_684 ();
 FILLCELL_X1 FILLER_114_688 ();
 FILLCELL_X32 FILLER_114_696 ();
 FILLCELL_X32 FILLER_114_728 ();
 FILLCELL_X2 FILLER_114_760 ();
 FILLCELL_X1 FILLER_114_766 ();
 FILLCELL_X4 FILLER_114_771 ();
 FILLCELL_X8 FILLER_114_778 ();
 FILLCELL_X4 FILLER_114_786 ();
 FILLCELL_X1 FILLER_114_790 ();
 FILLCELL_X4 FILLER_114_794 ();
 FILLCELL_X4 FILLER_114_805 ();
 FILLCELL_X4 FILLER_114_813 ();
 FILLCELL_X4 FILLER_114_830 ();
 FILLCELL_X1 FILLER_114_834 ();
 FILLCELL_X2 FILLER_114_845 ();
 FILLCELL_X1 FILLER_114_847 ();
 FILLCELL_X1 FILLER_114_856 ();
 FILLCELL_X1 FILLER_114_860 ();
 FILLCELL_X1 FILLER_114_876 ();
 FILLCELL_X2 FILLER_114_884 ();
 FILLCELL_X8 FILLER_114_902 ();
 FILLCELL_X1 FILLER_114_915 ();
 FILLCELL_X8 FILLER_114_941 ();
 FILLCELL_X16 FILLER_114_971 ();
 FILLCELL_X8 FILLER_114_987 ();
 FILLCELL_X4 FILLER_114_995 ();
 FILLCELL_X2 FILLER_114_999 ();
 FILLCELL_X1 FILLER_114_1016 ();
 FILLCELL_X1 FILLER_114_1028 ();
 FILLCELL_X1 FILLER_114_1040 ();
 FILLCELL_X1 FILLER_114_1050 ();
 FILLCELL_X2 FILLER_114_1063 ();
 FILLCELL_X2 FILLER_114_1103 ();
 FILLCELL_X1 FILLER_114_1105 ();
 FILLCELL_X2 FILLER_114_1119 ();
 FILLCELL_X1 FILLER_114_1121 ();
 FILLCELL_X4 FILLER_114_1126 ();
 FILLCELL_X2 FILLER_114_1146 ();
 FILLCELL_X8 FILLER_114_1154 ();
 FILLCELL_X2 FILLER_114_1173 ();
 FILLCELL_X16 FILLER_114_1187 ();
 FILLCELL_X4 FILLER_114_1203 ();
 FILLCELL_X2 FILLER_114_1207 ();
 FILLCELL_X32 FILLER_115_1 ();
 FILLCELL_X32 FILLER_115_33 ();
 FILLCELL_X32 FILLER_115_65 ();
 FILLCELL_X8 FILLER_115_97 ();
 FILLCELL_X4 FILLER_115_105 ();
 FILLCELL_X2 FILLER_115_109 ();
 FILLCELL_X1 FILLER_115_111 ();
 FILLCELL_X2 FILLER_115_129 ();
 FILLCELL_X8 FILLER_115_146 ();
 FILLCELL_X8 FILLER_115_158 ();
 FILLCELL_X4 FILLER_115_166 ();
 FILLCELL_X2 FILLER_115_182 ();
 FILLCELL_X1 FILLER_115_202 ();
 FILLCELL_X1 FILLER_115_209 ();
 FILLCELL_X2 FILLER_115_217 ();
 FILLCELL_X1 FILLER_115_219 ();
 FILLCELL_X2 FILLER_115_241 ();
 FILLCELL_X1 FILLER_115_248 ();
 FILLCELL_X2 FILLER_115_253 ();
 FILLCELL_X16 FILLER_115_286 ();
 FILLCELL_X4 FILLER_115_302 ();
 FILLCELL_X2 FILLER_115_310 ();
 FILLCELL_X2 FILLER_115_345 ();
 FILLCELL_X2 FILLER_115_357 ();
 FILLCELL_X1 FILLER_115_359 ();
 FILLCELL_X1 FILLER_115_374 ();
 FILLCELL_X2 FILLER_115_386 ();
 FILLCELL_X2 FILLER_115_392 ();
 FILLCELL_X2 FILLER_115_400 ();
 FILLCELL_X1 FILLER_115_402 ();
 FILLCELL_X4 FILLER_115_412 ();
 FILLCELL_X2 FILLER_115_419 ();
 FILLCELL_X1 FILLER_115_421 ();
 FILLCELL_X1 FILLER_115_426 ();
 FILLCELL_X8 FILLER_115_436 ();
 FILLCELL_X1 FILLER_115_444 ();
 FILLCELL_X1 FILLER_115_448 ();
 FILLCELL_X4 FILLER_115_459 ();
 FILLCELL_X32 FILLER_115_470 ();
 FILLCELL_X8 FILLER_115_502 ();
 FILLCELL_X4 FILLER_115_510 ();
 FILLCELL_X1 FILLER_115_514 ();
 FILLCELL_X1 FILLER_115_528 ();
 FILLCELL_X4 FILLER_115_535 ();
 FILLCELL_X2 FILLER_115_539 ();
 FILLCELL_X1 FILLER_115_541 ();
 FILLCELL_X4 FILLER_115_549 ();
 FILLCELL_X4 FILLER_115_563 ();
 FILLCELL_X4 FILLER_115_578 ();
 FILLCELL_X2 FILLER_115_582 ();
 FILLCELL_X8 FILLER_115_588 ();
 FILLCELL_X2 FILLER_115_596 ();
 FILLCELL_X2 FILLER_115_637 ();
 FILLCELL_X1 FILLER_115_639 ();
 FILLCELL_X2 FILLER_115_649 ();
 FILLCELL_X4 FILLER_115_658 ();
 FILLCELL_X1 FILLER_115_662 ();
 FILLCELL_X4 FILLER_115_676 ();
 FILLCELL_X2 FILLER_115_680 ();
 FILLCELL_X32 FILLER_115_713 ();
 FILLCELL_X16 FILLER_115_745 ();
 FILLCELL_X2 FILLER_115_765 ();
 FILLCELL_X2 FILLER_115_809 ();
 FILLCELL_X1 FILLER_115_811 ();
 FILLCELL_X16 FILLER_115_824 ();
 FILLCELL_X2 FILLER_115_840 ();
 FILLCELL_X1 FILLER_115_842 ();
 FILLCELL_X1 FILLER_115_861 ();
 FILLCELL_X8 FILLER_115_867 ();
 FILLCELL_X2 FILLER_115_875 ();
 FILLCELL_X1 FILLER_115_899 ();
 FILLCELL_X16 FILLER_115_903 ();
 FILLCELL_X2 FILLER_115_919 ();
 FILLCELL_X1 FILLER_115_938 ();
 FILLCELL_X4 FILLER_115_942 ();
 FILLCELL_X32 FILLER_115_960 ();
 FILLCELL_X8 FILLER_115_992 ();
 FILLCELL_X4 FILLER_115_1000 ();
 FILLCELL_X2 FILLER_115_1004 ();
 FILLCELL_X1 FILLER_115_1006 ();
 FILLCELL_X2 FILLER_115_1044 ();
 FILLCELL_X4 FILLER_115_1061 ();
 FILLCELL_X2 FILLER_115_1068 ();
 FILLCELL_X1 FILLER_115_1079 ();
 FILLCELL_X4 FILLER_115_1091 ();
 FILLCELL_X1 FILLER_115_1095 ();
 FILLCELL_X4 FILLER_115_1103 ();
 FILLCELL_X8 FILLER_115_1125 ();
 FILLCELL_X1 FILLER_115_1147 ();
 FILLCELL_X2 FILLER_115_1171 ();
 FILLCELL_X2 FILLER_115_1177 ();
 FILLCELL_X1 FILLER_115_1179 ();
 FILLCELL_X4 FILLER_115_1184 ();
 FILLCELL_X2 FILLER_115_1188 ();
 FILLCELL_X16 FILLER_115_1193 ();
 FILLCELL_X32 FILLER_116_1 ();
 FILLCELL_X32 FILLER_116_33 ();
 FILLCELL_X32 FILLER_116_65 ();
 FILLCELL_X4 FILLER_116_97 ();
 FILLCELL_X1 FILLER_116_101 ();
 FILLCELL_X1 FILLER_116_111 ();
 FILLCELL_X1 FILLER_116_120 ();
 FILLCELL_X1 FILLER_116_139 ();
 FILLCELL_X1 FILLER_116_144 ();
 FILLCELL_X1 FILLER_116_156 ();
 FILLCELL_X8 FILLER_116_161 ();
 FILLCELL_X4 FILLER_116_169 ();
 FILLCELL_X2 FILLER_116_173 ();
 FILLCELL_X1 FILLER_116_175 ();
 FILLCELL_X2 FILLER_116_195 ();
 FILLCELL_X1 FILLER_116_197 ();
 FILLCELL_X8 FILLER_116_214 ();
 FILLCELL_X2 FILLER_116_222 ();
 FILLCELL_X4 FILLER_116_227 ();
 FILLCELL_X8 FILLER_116_237 ();
 FILLCELL_X4 FILLER_116_245 ();
 FILLCELL_X2 FILLER_116_249 ();
 FILLCELL_X1 FILLER_116_251 ();
 FILLCELL_X32 FILLER_116_269 ();
 FILLCELL_X4 FILLER_116_301 ();
 FILLCELL_X1 FILLER_116_305 ();
 FILLCELL_X1 FILLER_116_313 ();
 FILLCELL_X2 FILLER_116_347 ();
 FILLCELL_X2 FILLER_116_354 ();
 FILLCELL_X2 FILLER_116_360 ();
 FILLCELL_X1 FILLER_116_385 ();
 FILLCELL_X2 FILLER_116_397 ();
 FILLCELL_X1 FILLER_116_399 ();
 FILLCELL_X1 FILLER_116_424 ();
 FILLCELL_X4 FILLER_116_428 ();
 FILLCELL_X2 FILLER_116_462 ();
 FILLCELL_X1 FILLER_116_464 ();
 FILLCELL_X32 FILLER_116_472 ();
 FILLCELL_X8 FILLER_116_504 ();
 FILLCELL_X4 FILLER_116_515 ();
 FILLCELL_X1 FILLER_116_519 ();
 FILLCELL_X4 FILLER_116_535 ();
 FILLCELL_X2 FILLER_116_539 ();
 FILLCELL_X1 FILLER_116_558 ();
 FILLCELL_X8 FILLER_116_574 ();
 FILLCELL_X16 FILLER_116_593 ();
 FILLCELL_X2 FILLER_116_609 ();
 FILLCELL_X1 FILLER_116_611 ();
 FILLCELL_X1 FILLER_116_619 ();
 FILLCELL_X1 FILLER_116_630 ();
 FILLCELL_X8 FILLER_116_645 ();
 FILLCELL_X1 FILLER_116_653 ();
 FILLCELL_X2 FILLER_116_675 ();
 FILLCELL_X16 FILLER_116_684 ();
 FILLCELL_X4 FILLER_116_700 ();
 FILLCELL_X2 FILLER_116_704 ();
 FILLCELL_X32 FILLER_116_709 ();
 FILLCELL_X16 FILLER_116_741 ();
 FILLCELL_X1 FILLER_116_757 ();
 FILLCELL_X4 FILLER_116_786 ();
 FILLCELL_X2 FILLER_116_790 ();
 FILLCELL_X1 FILLER_116_792 ();
 FILLCELL_X1 FILLER_116_798 ();
 FILLCELL_X4 FILLER_116_806 ();
 FILLCELL_X8 FILLER_116_813 ();
 FILLCELL_X1 FILLER_116_821 ();
 FILLCELL_X4 FILLER_116_827 ();
 FILLCELL_X2 FILLER_116_831 ();
 FILLCELL_X8 FILLER_116_837 ();
 FILLCELL_X4 FILLER_116_862 ();
 FILLCELL_X2 FILLER_116_870 ();
 FILLCELL_X1 FILLER_116_872 ();
 FILLCELL_X8 FILLER_116_878 ();
 FILLCELL_X2 FILLER_116_889 ();
 FILLCELL_X8 FILLER_116_909 ();
 FILLCELL_X1 FILLER_116_917 ();
 FILLCELL_X2 FILLER_116_925 ();
 FILLCELL_X1 FILLER_116_927 ();
 FILLCELL_X4 FILLER_116_933 ();
 FILLCELL_X4 FILLER_116_942 ();
 FILLCELL_X2 FILLER_116_946 ();
 FILLCELL_X1 FILLER_116_948 ();
 FILLCELL_X8 FILLER_116_962 ();
 FILLCELL_X4 FILLER_116_970 ();
 FILLCELL_X1 FILLER_116_974 ();
 FILLCELL_X4 FILLER_116_980 ();
 FILLCELL_X1 FILLER_116_984 ();
 FILLCELL_X2 FILLER_116_1027 ();
 FILLCELL_X2 FILLER_116_1074 ();
 FILLCELL_X4 FILLER_116_1079 ();
 FILLCELL_X4 FILLER_116_1090 ();
 FILLCELL_X1 FILLER_116_1108 ();
 FILLCELL_X4 FILLER_116_1112 ();
 FILLCELL_X2 FILLER_116_1128 ();
 FILLCELL_X1 FILLER_116_1130 ();
 FILLCELL_X1 FILLER_116_1146 ();
 FILLCELL_X1 FILLER_116_1151 ();
 FILLCELL_X2 FILLER_116_1157 ();
 FILLCELL_X1 FILLER_116_1159 ();
 FILLCELL_X1 FILLER_116_1166 ();
 FILLCELL_X2 FILLER_116_1171 ();
 FILLCELL_X1 FILLER_116_1173 ();
 FILLCELL_X16 FILLER_116_1184 ();
 FILLCELL_X8 FILLER_116_1200 ();
 FILLCELL_X1 FILLER_116_1208 ();
 FILLCELL_X32 FILLER_117_1 ();
 FILLCELL_X32 FILLER_117_33 ();
 FILLCELL_X32 FILLER_117_65 ();
 FILLCELL_X1 FILLER_117_97 ();
 FILLCELL_X4 FILLER_117_105 ();
 FILLCELL_X2 FILLER_117_109 ();
 FILLCELL_X2 FILLER_117_149 ();
 FILLCELL_X1 FILLER_117_160 ();
 FILLCELL_X2 FILLER_117_168 ();
 FILLCELL_X4 FILLER_117_173 ();
 FILLCELL_X2 FILLER_117_177 ();
 FILLCELL_X1 FILLER_117_184 ();
 FILLCELL_X2 FILLER_117_189 ();
 FILLCELL_X4 FILLER_117_202 ();
 FILLCELL_X1 FILLER_117_211 ();
 FILLCELL_X2 FILLER_117_221 ();
 FILLCELL_X2 FILLER_117_228 ();
 FILLCELL_X1 FILLER_117_260 ();
 FILLCELL_X16 FILLER_117_264 ();
 FILLCELL_X4 FILLER_117_280 ();
 FILLCELL_X1 FILLER_117_284 ();
 FILLCELL_X4 FILLER_117_319 ();
 FILLCELL_X2 FILLER_117_323 ();
 FILLCELL_X2 FILLER_117_333 ();
 FILLCELL_X4 FILLER_117_339 ();
 FILLCELL_X2 FILLER_117_343 ();
 FILLCELL_X2 FILLER_117_353 ();
 FILLCELL_X4 FILLER_117_362 ();
 FILLCELL_X8 FILLER_117_370 ();
 FILLCELL_X1 FILLER_117_378 ();
 FILLCELL_X2 FILLER_117_383 ();
 FILLCELL_X4 FILLER_117_394 ();
 FILLCELL_X2 FILLER_117_398 ();
 FILLCELL_X1 FILLER_117_400 ();
 FILLCELL_X8 FILLER_117_412 ();
 FILLCELL_X1 FILLER_117_420 ();
 FILLCELL_X1 FILLER_117_452 ();
 FILLCELL_X2 FILLER_117_457 ();
 FILLCELL_X32 FILLER_117_466 ();
 FILLCELL_X8 FILLER_117_498 ();
 FILLCELL_X4 FILLER_117_506 ();
 FILLCELL_X1 FILLER_117_510 ();
 FILLCELL_X4 FILLER_117_521 ();
 FILLCELL_X1 FILLER_117_525 ();
 FILLCELL_X1 FILLER_117_548 ();
 FILLCELL_X4 FILLER_117_563 ();
 FILLCELL_X1 FILLER_117_567 ();
 FILLCELL_X2 FILLER_117_598 ();
 FILLCELL_X4 FILLER_117_610 ();
 FILLCELL_X1 FILLER_117_624 ();
 FILLCELL_X8 FILLER_117_635 ();
 FILLCELL_X16 FILLER_117_669 ();
 FILLCELL_X8 FILLER_117_685 ();
 FILLCELL_X2 FILLER_117_693 ();
 FILLCELL_X1 FILLER_117_695 ();
 FILLCELL_X2 FILLER_117_717 ();
 FILLCELL_X1 FILLER_117_719 ();
 FILLCELL_X16 FILLER_117_727 ();
 FILLCELL_X8 FILLER_117_743 ();
 FILLCELL_X4 FILLER_117_751 ();
 FILLCELL_X2 FILLER_117_755 ();
 FILLCELL_X8 FILLER_117_771 ();
 FILLCELL_X1 FILLER_117_783 ();
 FILLCELL_X2 FILLER_117_797 ();
 FILLCELL_X1 FILLER_117_799 ();
 FILLCELL_X1 FILLER_117_815 ();
 FILLCELL_X1 FILLER_117_818 ();
 FILLCELL_X1 FILLER_117_831 ();
 FILLCELL_X4 FILLER_117_837 ();
 FILLCELL_X2 FILLER_117_856 ();
 FILLCELL_X1 FILLER_117_871 ();
 FILLCELL_X2 FILLER_117_888 ();
 FILLCELL_X2 FILLER_117_897 ();
 FILLCELL_X8 FILLER_117_912 ();
 FILLCELL_X1 FILLER_117_930 ();
 FILLCELL_X8 FILLER_117_938 ();
 FILLCELL_X1 FILLER_117_946 ();
 FILLCELL_X16 FILLER_117_960 ();
 FILLCELL_X4 FILLER_117_976 ();
 FILLCELL_X2 FILLER_117_980 ();
 FILLCELL_X1 FILLER_117_982 ();
 FILLCELL_X8 FILLER_117_988 ();
 FILLCELL_X2 FILLER_117_996 ();
 FILLCELL_X1 FILLER_117_998 ();
 FILLCELL_X2 FILLER_117_1016 ();
 FILLCELL_X1 FILLER_117_1018 ();
 FILLCELL_X2 FILLER_117_1091 ();
 FILLCELL_X2 FILLER_117_1114 ();
 FILLCELL_X1 FILLER_117_1116 ();
 FILLCELL_X8 FILLER_117_1121 ();
 FILLCELL_X4 FILLER_117_1129 ();
 FILLCELL_X4 FILLER_117_1138 ();
 FILLCELL_X2 FILLER_117_1142 ();
 FILLCELL_X1 FILLER_117_1144 ();
 FILLCELL_X16 FILLER_117_1149 ();
 FILLCELL_X2 FILLER_117_1174 ();
 FILLCELL_X1 FILLER_117_1176 ();
 FILLCELL_X16 FILLER_117_1182 ();
 FILLCELL_X8 FILLER_117_1198 ();
 FILLCELL_X2 FILLER_117_1206 ();
 FILLCELL_X1 FILLER_117_1208 ();
 FILLCELL_X32 FILLER_118_1 ();
 FILLCELL_X32 FILLER_118_33 ();
 FILLCELL_X32 FILLER_118_65 ();
 FILLCELL_X4 FILLER_118_97 ();
 FILLCELL_X1 FILLER_118_101 ();
 FILLCELL_X1 FILLER_118_161 ();
 FILLCELL_X1 FILLER_118_166 ();
 FILLCELL_X8 FILLER_118_178 ();
 FILLCELL_X2 FILLER_118_204 ();
 FILLCELL_X1 FILLER_118_223 ();
 FILLCELL_X2 FILLER_118_242 ();
 FILLCELL_X1 FILLER_118_244 ();
 FILLCELL_X16 FILLER_118_267 ();
 FILLCELL_X8 FILLER_118_283 ();
 FILLCELL_X2 FILLER_118_305 ();
 FILLCELL_X2 FILLER_118_316 ();
 FILLCELL_X1 FILLER_118_318 ();
 FILLCELL_X2 FILLER_118_323 ();
 FILLCELL_X2 FILLER_118_331 ();
 FILLCELL_X4 FILLER_118_344 ();
 FILLCELL_X1 FILLER_118_348 ();
 FILLCELL_X4 FILLER_118_353 ();
 FILLCELL_X1 FILLER_118_357 ();
 FILLCELL_X2 FILLER_118_371 ();
 FILLCELL_X16 FILLER_118_381 ();
 FILLCELL_X8 FILLER_118_397 ();
 FILLCELL_X1 FILLER_118_405 ();
 FILLCELL_X1 FILLER_118_415 ();
 FILLCELL_X2 FILLER_118_422 ();
 FILLCELL_X1 FILLER_118_436 ();
 FILLCELL_X2 FILLER_118_446 ();
 FILLCELL_X2 FILLER_118_455 ();
 FILLCELL_X1 FILLER_118_457 ();
 FILLCELL_X1 FILLER_118_469 ();
 FILLCELL_X8 FILLER_118_484 ();
 FILLCELL_X1 FILLER_118_492 ();
 FILLCELL_X16 FILLER_118_515 ();
 FILLCELL_X8 FILLER_118_541 ();
 FILLCELL_X1 FILLER_118_549 ();
 FILLCELL_X16 FILLER_118_560 ();
 FILLCELL_X1 FILLER_118_576 ();
 FILLCELL_X8 FILLER_118_591 ();
 FILLCELL_X16 FILLER_118_606 ();
 FILLCELL_X8 FILLER_118_622 ();
 FILLCELL_X1 FILLER_118_630 ();
 FILLCELL_X2 FILLER_118_632 ();
 FILLCELL_X1 FILLER_118_634 ();
 FILLCELL_X8 FILLER_118_684 ();
 FILLCELL_X4 FILLER_118_692 ();
 FILLCELL_X2 FILLER_118_696 ();
 FILLCELL_X8 FILLER_118_705 ();
 FILLCELL_X2 FILLER_118_713 ();
 FILLCELL_X2 FILLER_118_721 ();
 FILLCELL_X8 FILLER_118_747 ();
 FILLCELL_X2 FILLER_118_755 ();
 FILLCELL_X2 FILLER_118_761 ();
 FILLCELL_X1 FILLER_118_763 ();
 FILLCELL_X1 FILLER_118_772 ();
 FILLCELL_X2 FILLER_118_777 ();
 FILLCELL_X8 FILLER_118_795 ();
 FILLCELL_X4 FILLER_118_809 ();
 FILLCELL_X1 FILLER_118_813 ();
 FILLCELL_X2 FILLER_118_822 ();
 FILLCELL_X1 FILLER_118_839 ();
 FILLCELL_X2 FILLER_118_851 ();
 FILLCELL_X8 FILLER_118_869 ();
 FILLCELL_X2 FILLER_118_887 ();
 FILLCELL_X2 FILLER_118_896 ();
 FILLCELL_X4 FILLER_118_914 ();
 FILLCELL_X1 FILLER_118_929 ();
 FILLCELL_X2 FILLER_118_941 ();
 FILLCELL_X32 FILLER_118_960 ();
 FILLCELL_X16 FILLER_118_992 ();
 FILLCELL_X8 FILLER_118_1008 ();
 FILLCELL_X1 FILLER_118_1016 ();
 FILLCELL_X1 FILLER_118_1030 ();
 FILLCELL_X1 FILLER_118_1076 ();
 FILLCELL_X2 FILLER_118_1083 ();
 FILLCELL_X1 FILLER_118_1099 ();
 FILLCELL_X2 FILLER_118_1114 ();
 FILLCELL_X1 FILLER_118_1116 ();
 FILLCELL_X1 FILLER_118_1125 ();
 FILLCELL_X1 FILLER_118_1129 ();
 FILLCELL_X2 FILLER_118_1141 ();
 FILLCELL_X4 FILLER_118_1147 ();
 FILLCELL_X4 FILLER_118_1161 ();
 FILLCELL_X1 FILLER_118_1165 ();
 FILLCELL_X32 FILLER_118_1170 ();
 FILLCELL_X4 FILLER_118_1202 ();
 FILLCELL_X2 FILLER_118_1206 ();
 FILLCELL_X1 FILLER_118_1208 ();
 FILLCELL_X32 FILLER_119_1 ();
 FILLCELL_X32 FILLER_119_33 ();
 FILLCELL_X32 FILLER_119_65 ();
 FILLCELL_X4 FILLER_119_97 ();
 FILLCELL_X1 FILLER_119_101 ();
 FILLCELL_X2 FILLER_119_109 ();
 FILLCELL_X1 FILLER_119_120 ();
 FILLCELL_X2 FILLER_119_132 ();
 FILLCELL_X2 FILLER_119_152 ();
 FILLCELL_X1 FILLER_119_189 ();
 FILLCELL_X1 FILLER_119_193 ();
 FILLCELL_X1 FILLER_119_205 ();
 FILLCELL_X1 FILLER_119_210 ();
 FILLCELL_X2 FILLER_119_221 ();
 FILLCELL_X1 FILLER_119_223 ();
 FILLCELL_X4 FILLER_119_233 ();
 FILLCELL_X2 FILLER_119_237 ();
 FILLCELL_X1 FILLER_119_239 ();
 FILLCELL_X4 FILLER_119_245 ();
 FILLCELL_X1 FILLER_119_249 ();
 FILLCELL_X16 FILLER_119_263 ();
 FILLCELL_X8 FILLER_119_279 ();
 FILLCELL_X1 FILLER_119_312 ();
 FILLCELL_X2 FILLER_119_316 ();
 FILLCELL_X4 FILLER_119_324 ();
 FILLCELL_X8 FILLER_119_335 ();
 FILLCELL_X4 FILLER_119_343 ();
 FILLCELL_X1 FILLER_119_347 ();
 FILLCELL_X4 FILLER_119_357 ();
 FILLCELL_X2 FILLER_119_402 ();
 FILLCELL_X1 FILLER_119_414 ();
 FILLCELL_X2 FILLER_119_426 ();
 FILLCELL_X1 FILLER_119_428 ();
 FILLCELL_X2 FILLER_119_433 ();
 FILLCELL_X1 FILLER_119_438 ();
 FILLCELL_X1 FILLER_119_447 ();
 FILLCELL_X2 FILLER_119_466 ();
 FILLCELL_X1 FILLER_119_468 ();
 FILLCELL_X16 FILLER_119_482 ();
 FILLCELL_X8 FILLER_119_498 ();
 FILLCELL_X2 FILLER_119_506 ();
 FILLCELL_X32 FILLER_119_514 ();
 FILLCELL_X8 FILLER_119_546 ();
 FILLCELL_X4 FILLER_119_554 ();
 FILLCELL_X2 FILLER_119_558 ();
 FILLCELL_X16 FILLER_119_586 ();
 FILLCELL_X2 FILLER_119_602 ();
 FILLCELL_X1 FILLER_119_604 ();
 FILLCELL_X32 FILLER_119_611 ();
 FILLCELL_X16 FILLER_119_643 ();
 FILLCELL_X2 FILLER_119_659 ();
 FILLCELL_X1 FILLER_119_661 ();
 FILLCELL_X8 FILLER_119_694 ();
 FILLCELL_X2 FILLER_119_702 ();
 FILLCELL_X1 FILLER_119_704 ();
 FILLCELL_X1 FILLER_119_734 ();
 FILLCELL_X16 FILLER_119_740 ();
 FILLCELL_X2 FILLER_119_756 ();
 FILLCELL_X1 FILLER_119_758 ();
 FILLCELL_X1 FILLER_119_763 ();
 FILLCELL_X1 FILLER_119_767 ();
 FILLCELL_X4 FILLER_119_797 ();
 FILLCELL_X2 FILLER_119_801 ();
 FILLCELL_X1 FILLER_119_803 ();
 FILLCELL_X4 FILLER_119_808 ();
 FILLCELL_X2 FILLER_119_812 ();
 FILLCELL_X4 FILLER_119_825 ();
 FILLCELL_X2 FILLER_119_837 ();
 FILLCELL_X4 FILLER_119_852 ();
 FILLCELL_X4 FILLER_119_862 ();
 FILLCELL_X1 FILLER_119_880 ();
 FILLCELL_X2 FILLER_119_885 ();
 FILLCELL_X1 FILLER_119_899 ();
 FILLCELL_X2 FILLER_119_904 ();
 FILLCELL_X8 FILLER_119_914 ();
 FILLCELL_X1 FILLER_119_922 ();
 FILLCELL_X8 FILLER_119_934 ();
 FILLCELL_X4 FILLER_119_942 ();
 FILLCELL_X2 FILLER_119_946 ();
 FILLCELL_X16 FILLER_119_962 ();
 FILLCELL_X2 FILLER_119_978 ();
 FILLCELL_X16 FILLER_119_993 ();
 FILLCELL_X1 FILLER_119_1009 ();
 FILLCELL_X2 FILLER_119_1080 ();
 FILLCELL_X16 FILLER_119_1092 ();
 FILLCELL_X8 FILLER_119_1108 ();
 FILLCELL_X2 FILLER_119_1116 ();
 FILLCELL_X1 FILLER_119_1123 ();
 FILLCELL_X2 FILLER_119_1127 ();
 FILLCELL_X2 FILLER_119_1147 ();
 FILLCELL_X4 FILLER_119_1161 ();
 FILLCELL_X16 FILLER_119_1185 ();
 FILLCELL_X8 FILLER_119_1201 ();
 FILLCELL_X32 FILLER_120_1 ();
 FILLCELL_X32 FILLER_120_33 ();
 FILLCELL_X32 FILLER_120_65 ();
 FILLCELL_X8 FILLER_120_97 ();
 FILLCELL_X2 FILLER_120_105 ();
 FILLCELL_X1 FILLER_120_107 ();
 FILLCELL_X4 FILLER_120_161 ();
 FILLCELL_X1 FILLER_120_172 ();
 FILLCELL_X1 FILLER_120_180 ();
 FILLCELL_X4 FILLER_120_210 ();
 FILLCELL_X2 FILLER_120_214 ();
 FILLCELL_X1 FILLER_120_216 ();
 FILLCELL_X8 FILLER_120_224 ();
 FILLCELL_X4 FILLER_120_236 ();
 FILLCELL_X1 FILLER_120_260 ();
 FILLCELL_X16 FILLER_120_265 ();
 FILLCELL_X8 FILLER_120_281 ();
 FILLCELL_X4 FILLER_120_289 ();
 FILLCELL_X2 FILLER_120_293 ();
 FILLCELL_X1 FILLER_120_295 ();
 FILLCELL_X2 FILLER_120_376 ();
 FILLCELL_X2 FILLER_120_397 ();
 FILLCELL_X1 FILLER_120_399 ();
 FILLCELL_X4 FILLER_120_422 ();
 FILLCELL_X2 FILLER_120_426 ();
 FILLCELL_X1 FILLER_120_428 ();
 FILLCELL_X2 FILLER_120_437 ();
 FILLCELL_X4 FILLER_120_444 ();
 FILLCELL_X1 FILLER_120_448 ();
 FILLCELL_X32 FILLER_120_453 ();
 FILLCELL_X16 FILLER_120_485 ();
 FILLCELL_X8 FILLER_120_501 ();
 FILLCELL_X1 FILLER_120_509 ();
 FILLCELL_X1 FILLER_120_517 ();
 FILLCELL_X16 FILLER_120_545 ();
 FILLCELL_X2 FILLER_120_561 ();
 FILLCELL_X1 FILLER_120_563 ();
 FILLCELL_X4 FILLER_120_605 ();
 FILLCELL_X4 FILLER_120_626 ();
 FILLCELL_X1 FILLER_120_630 ();
 FILLCELL_X4 FILLER_120_632 ();
 FILLCELL_X2 FILLER_120_636 ();
 FILLCELL_X2 FILLER_120_642 ();
 FILLCELL_X1 FILLER_120_652 ();
 FILLCELL_X2 FILLER_120_656 ();
 FILLCELL_X1 FILLER_120_658 ();
 FILLCELL_X4 FILLER_120_683 ();
 FILLCELL_X1 FILLER_120_687 ();
 FILLCELL_X2 FILLER_120_705 ();
 FILLCELL_X16 FILLER_120_737 ();
 FILLCELL_X4 FILLER_120_753 ();
 FILLCELL_X2 FILLER_120_757 ();
 FILLCELL_X2 FILLER_120_777 ();
 FILLCELL_X1 FILLER_120_779 ();
 FILLCELL_X8 FILLER_120_793 ();
 FILLCELL_X1 FILLER_120_801 ();
 FILLCELL_X8 FILLER_120_812 ();
 FILLCELL_X2 FILLER_120_820 ();
 FILLCELL_X1 FILLER_120_822 ();
 FILLCELL_X4 FILLER_120_827 ();
 FILLCELL_X2 FILLER_120_831 ();
 FILLCELL_X4 FILLER_120_837 ();
 FILLCELL_X2 FILLER_120_841 ();
 FILLCELL_X4 FILLER_120_846 ();
 FILLCELL_X1 FILLER_120_850 ();
 FILLCELL_X2 FILLER_120_859 ();
 FILLCELL_X1 FILLER_120_872 ();
 FILLCELL_X4 FILLER_120_902 ();
 FILLCELL_X2 FILLER_120_906 ();
 FILLCELL_X1 FILLER_120_928 ();
 FILLCELL_X4 FILLER_120_951 ();
 FILLCELL_X2 FILLER_120_955 ();
 FILLCELL_X1 FILLER_120_957 ();
 FILLCELL_X16 FILLER_120_962 ();
 FILLCELL_X8 FILLER_120_978 ();
 FILLCELL_X2 FILLER_120_986 ();
 FILLCELL_X1 FILLER_120_988 ();
 FILLCELL_X8 FILLER_120_1013 ();
 FILLCELL_X1 FILLER_120_1021 ();
 FILLCELL_X2 FILLER_120_1034 ();
 FILLCELL_X1 FILLER_120_1036 ();
 FILLCELL_X2 FILLER_120_1067 ();
 FILLCELL_X1 FILLER_120_1069 ();
 FILLCELL_X2 FILLER_120_1077 ();
 FILLCELL_X2 FILLER_120_1086 ();
 FILLCELL_X1 FILLER_120_1097 ();
 FILLCELL_X1 FILLER_120_1127 ();
 FILLCELL_X1 FILLER_120_1133 ();
 FILLCELL_X2 FILLER_120_1147 ();
 FILLCELL_X32 FILLER_120_1170 ();
 FILLCELL_X4 FILLER_120_1202 ();
 FILLCELL_X2 FILLER_120_1206 ();
 FILLCELL_X1 FILLER_120_1208 ();
 FILLCELL_X32 FILLER_121_1 ();
 FILLCELL_X32 FILLER_121_33 ();
 FILLCELL_X32 FILLER_121_65 ();
 FILLCELL_X16 FILLER_121_97 ();
 FILLCELL_X4 FILLER_121_113 ();
 FILLCELL_X1 FILLER_121_135 ();
 FILLCELL_X1 FILLER_121_162 ();
 FILLCELL_X1 FILLER_121_166 ();
 FILLCELL_X2 FILLER_121_193 ();
 FILLCELL_X1 FILLER_121_223 ();
 FILLCELL_X16 FILLER_121_262 ();
 FILLCELL_X8 FILLER_121_278 ();
 FILLCELL_X4 FILLER_121_286 ();
 FILLCELL_X1 FILLER_121_290 ();
 FILLCELL_X4 FILLER_121_302 ();
 FILLCELL_X1 FILLER_121_306 ();
 FILLCELL_X1 FILLER_121_311 ();
 FILLCELL_X1 FILLER_121_316 ();
 FILLCELL_X2 FILLER_121_325 ();
 FILLCELL_X4 FILLER_121_352 ();
 FILLCELL_X1 FILLER_121_356 ();
 FILLCELL_X4 FILLER_121_360 ();
 FILLCELL_X2 FILLER_121_364 ();
 FILLCELL_X1 FILLER_121_366 ();
 FILLCELL_X4 FILLER_121_376 ();
 FILLCELL_X2 FILLER_121_380 ();
 FILLCELL_X2 FILLER_121_400 ();
 FILLCELL_X1 FILLER_121_402 ();
 FILLCELL_X2 FILLER_121_408 ();
 FILLCELL_X2 FILLER_121_414 ();
 FILLCELL_X1 FILLER_121_431 ();
 FILLCELL_X2 FILLER_121_437 ();
 FILLCELL_X1 FILLER_121_439 ();
 FILLCELL_X8 FILLER_121_481 ();
 FILLCELL_X2 FILLER_121_489 ();
 FILLCELL_X1 FILLER_121_491 ();
 FILLCELL_X4 FILLER_121_519 ();
 FILLCELL_X2 FILLER_121_523 ();
 FILLCELL_X4 FILLER_121_559 ();
 FILLCELL_X2 FILLER_121_599 ();
 FILLCELL_X2 FILLER_121_634 ();
 FILLCELL_X8 FILLER_121_660 ();
 FILLCELL_X4 FILLER_121_668 ();
 FILLCELL_X16 FILLER_121_680 ();
 FILLCELL_X8 FILLER_121_696 ();
 FILLCELL_X2 FILLER_121_704 ();
 FILLCELL_X32 FILLER_121_716 ();
 FILLCELL_X1 FILLER_121_759 ();
 FILLCELL_X1 FILLER_121_768 ();
 FILLCELL_X1 FILLER_121_773 ();
 FILLCELL_X2 FILLER_121_778 ();
 FILLCELL_X1 FILLER_121_780 ();
 FILLCELL_X2 FILLER_121_785 ();
 FILLCELL_X1 FILLER_121_787 ();
 FILLCELL_X8 FILLER_121_791 ();
 FILLCELL_X32 FILLER_121_802 ();
 FILLCELL_X1 FILLER_121_834 ();
 FILLCELL_X1 FILLER_121_865 ();
 FILLCELL_X2 FILLER_121_870 ();
 FILLCELL_X1 FILLER_121_872 ();
 FILLCELL_X2 FILLER_121_878 ();
 FILLCELL_X4 FILLER_121_909 ();
 FILLCELL_X1 FILLER_121_937 ();
 FILLCELL_X1 FILLER_121_955 ();
 FILLCELL_X16 FILLER_121_978 ();
 FILLCELL_X2 FILLER_121_994 ();
 FILLCELL_X1 FILLER_121_996 ();
 FILLCELL_X2 FILLER_121_1006 ();
 FILLCELL_X2 FILLER_121_1056 ();
 FILLCELL_X1 FILLER_121_1058 ();
 FILLCELL_X4 FILLER_121_1122 ();
 FILLCELL_X2 FILLER_121_1126 ();
 FILLCELL_X4 FILLER_121_1138 ();
 FILLCELL_X2 FILLER_121_1142 ();
 FILLCELL_X16 FILLER_121_1193 ();
 FILLCELL_X32 FILLER_122_1 ();
 FILLCELL_X32 FILLER_122_33 ();
 FILLCELL_X32 FILLER_122_65 ();
 FILLCELL_X16 FILLER_122_97 ();
 FILLCELL_X8 FILLER_122_113 ();
 FILLCELL_X2 FILLER_122_121 ();
 FILLCELL_X1 FILLER_122_123 ();
 FILLCELL_X1 FILLER_122_135 ();
 FILLCELL_X2 FILLER_122_158 ();
 FILLCELL_X4 FILLER_122_170 ();
 FILLCELL_X1 FILLER_122_174 ();
 FILLCELL_X2 FILLER_122_186 ();
 FILLCELL_X1 FILLER_122_188 ();
 FILLCELL_X2 FILLER_122_202 ();
 FILLCELL_X8 FILLER_122_218 ();
 FILLCELL_X1 FILLER_122_226 ();
 FILLCELL_X32 FILLER_122_249 ();
 FILLCELL_X2 FILLER_122_281 ();
 FILLCELL_X1 FILLER_122_283 ();
 FILLCELL_X1 FILLER_122_294 ();
 FILLCELL_X2 FILLER_122_299 ();
 FILLCELL_X2 FILLER_122_314 ();
 FILLCELL_X2 FILLER_122_320 ();
 FILLCELL_X1 FILLER_122_322 ();
 FILLCELL_X4 FILLER_122_329 ();
 FILLCELL_X4 FILLER_122_369 ();
 FILLCELL_X1 FILLER_122_373 ();
 FILLCELL_X8 FILLER_122_415 ();
 FILLCELL_X4 FILLER_122_423 ();
 FILLCELL_X2 FILLER_122_427 ();
 FILLCELL_X1 FILLER_122_429 ();
 FILLCELL_X8 FILLER_122_434 ();
 FILLCELL_X4 FILLER_122_442 ();
 FILLCELL_X1 FILLER_122_446 ();
 FILLCELL_X4 FILLER_122_455 ();
 FILLCELL_X32 FILLER_122_466 ();
 FILLCELL_X2 FILLER_122_498 ();
 FILLCELL_X1 FILLER_122_500 ();
 FILLCELL_X4 FILLER_122_504 ();
 FILLCELL_X2 FILLER_122_539 ();
 FILLCELL_X8 FILLER_122_569 ();
 FILLCELL_X1 FILLER_122_577 ();
 FILLCELL_X8 FILLER_122_596 ();
 FILLCELL_X2 FILLER_122_620 ();
 FILLCELL_X2 FILLER_122_629 ();
 FILLCELL_X2 FILLER_122_632 ();
 FILLCELL_X1 FILLER_122_634 ();
 FILLCELL_X4 FILLER_122_698 ();
 FILLCELL_X1 FILLER_122_702 ();
 FILLCELL_X4 FILLER_122_710 ();
 FILLCELL_X2 FILLER_122_714 ();
 FILLCELL_X1 FILLER_122_716 ();
 FILLCELL_X16 FILLER_122_734 ();
 FILLCELL_X4 FILLER_122_750 ();
 FILLCELL_X2 FILLER_122_754 ();
 FILLCELL_X1 FILLER_122_756 ();
 FILLCELL_X2 FILLER_122_768 ();
 FILLCELL_X1 FILLER_122_779 ();
 FILLCELL_X8 FILLER_122_792 ();
 FILLCELL_X1 FILLER_122_800 ();
 FILLCELL_X4 FILLER_122_804 ();
 FILLCELL_X1 FILLER_122_808 ();
 FILLCELL_X32 FILLER_122_817 ();
 FILLCELL_X4 FILLER_122_849 ();
 FILLCELL_X2 FILLER_122_853 ();
 FILLCELL_X1 FILLER_122_855 ();
 FILLCELL_X8 FILLER_122_864 ();
 FILLCELL_X2 FILLER_122_872 ();
 FILLCELL_X1 FILLER_122_887 ();
 FILLCELL_X8 FILLER_122_895 ();
 FILLCELL_X4 FILLER_122_905 ();
 FILLCELL_X2 FILLER_122_909 ();
 FILLCELL_X1 FILLER_122_911 ();
 FILLCELL_X2 FILLER_122_916 ();
 FILLCELL_X1 FILLER_122_926 ();
 FILLCELL_X8 FILLER_122_959 ();
 FILLCELL_X4 FILLER_122_967 ();
 FILLCELL_X2 FILLER_122_971 ();
 FILLCELL_X1 FILLER_122_973 ();
 FILLCELL_X16 FILLER_122_980 ();
 FILLCELL_X2 FILLER_122_1006 ();
 FILLCELL_X1 FILLER_122_1008 ();
 FILLCELL_X32 FILLER_122_1026 ();
 FILLCELL_X8 FILLER_122_1058 ();
 FILLCELL_X4 FILLER_122_1066 ();
 FILLCELL_X2 FILLER_122_1070 ();
 FILLCELL_X16 FILLER_122_1076 ();
 FILLCELL_X8 FILLER_122_1092 ();
 FILLCELL_X2 FILLER_122_1100 ();
 FILLCELL_X1 FILLER_122_1102 ();
 FILLCELL_X2 FILLER_122_1113 ();
 FILLCELL_X32 FILLER_122_1132 ();
 FILLCELL_X32 FILLER_122_1164 ();
 FILLCELL_X8 FILLER_122_1196 ();
 FILLCELL_X4 FILLER_122_1204 ();
 FILLCELL_X1 FILLER_122_1208 ();
 FILLCELL_X32 FILLER_123_1 ();
 FILLCELL_X32 FILLER_123_33 ();
 FILLCELL_X32 FILLER_123_65 ();
 FILLCELL_X16 FILLER_123_97 ();
 FILLCELL_X2 FILLER_123_113 ();
 FILLCELL_X4 FILLER_123_130 ();
 FILLCELL_X2 FILLER_123_150 ();
 FILLCELL_X1 FILLER_123_152 ();
 FILLCELL_X2 FILLER_123_158 ();
 FILLCELL_X2 FILLER_123_225 ();
 FILLCELL_X2 FILLER_123_232 ();
 FILLCELL_X2 FILLER_123_237 ();
 FILLCELL_X2 FILLER_123_244 ();
 FILLCELL_X16 FILLER_123_262 ();
 FILLCELL_X2 FILLER_123_278 ();
 FILLCELL_X1 FILLER_123_280 ();
 FILLCELL_X2 FILLER_123_323 ();
 FILLCELL_X1 FILLER_123_325 ();
 FILLCELL_X8 FILLER_123_333 ();
 FILLCELL_X1 FILLER_123_341 ();
 FILLCELL_X1 FILLER_123_365 ();
 FILLCELL_X1 FILLER_123_369 ();
 FILLCELL_X2 FILLER_123_374 ();
 FILLCELL_X2 FILLER_123_387 ();
 FILLCELL_X1 FILLER_123_393 ();
 FILLCELL_X1 FILLER_123_401 ();
 FILLCELL_X8 FILLER_123_413 ();
 FILLCELL_X4 FILLER_123_421 ();
 FILLCELL_X4 FILLER_123_437 ();
 FILLCELL_X1 FILLER_123_441 ();
 FILLCELL_X4 FILLER_123_446 ();
 FILLCELL_X2 FILLER_123_455 ();
 FILLCELL_X1 FILLER_123_457 ();
 FILLCELL_X32 FILLER_123_463 ();
 FILLCELL_X16 FILLER_123_495 ();
 FILLCELL_X8 FILLER_123_511 ();
 FILLCELL_X1 FILLER_123_519 ();
 FILLCELL_X1 FILLER_123_533 ();
 FILLCELL_X8 FILLER_123_565 ();
 FILLCELL_X2 FILLER_123_573 ();
 FILLCELL_X1 FILLER_123_575 ();
 FILLCELL_X4 FILLER_123_585 ();
 FILLCELL_X2 FILLER_123_589 ();
 FILLCELL_X1 FILLER_123_591 ();
 FILLCELL_X2 FILLER_123_595 ();
 FILLCELL_X2 FILLER_123_600 ();
 FILLCELL_X2 FILLER_123_608 ();
 FILLCELL_X1 FILLER_123_610 ();
 FILLCELL_X2 FILLER_123_621 ();
 FILLCELL_X16 FILLER_123_647 ();
 FILLCELL_X2 FILLER_123_670 ();
 FILLCELL_X1 FILLER_123_678 ();
 FILLCELL_X4 FILLER_123_696 ();
 FILLCELL_X2 FILLER_123_700 ();
 FILLCELL_X8 FILLER_123_716 ();
 FILLCELL_X8 FILLER_123_741 ();
 FILLCELL_X4 FILLER_123_749 ();
 FILLCELL_X2 FILLER_123_775 ();
 FILLCELL_X1 FILLER_123_777 ();
 FILLCELL_X8 FILLER_123_799 ();
 FILLCELL_X2 FILLER_123_818 ();
 FILLCELL_X1 FILLER_123_826 ();
 FILLCELL_X4 FILLER_123_835 ();
 FILLCELL_X1 FILLER_123_839 ();
 FILLCELL_X1 FILLER_123_845 ();
 FILLCELL_X4 FILLER_123_869 ();
 FILLCELL_X2 FILLER_123_873 ();
 FILLCELL_X1 FILLER_123_875 ();
 FILLCELL_X8 FILLER_123_883 ();
 FILLCELL_X2 FILLER_123_891 ();
 FILLCELL_X1 FILLER_123_893 ();
 FILLCELL_X2 FILLER_123_902 ();
 FILLCELL_X1 FILLER_123_944 ();
 FILLCELL_X1 FILLER_123_958 ();
 FILLCELL_X8 FILLER_123_966 ();
 FILLCELL_X8 FILLER_123_980 ();
 FILLCELL_X4 FILLER_123_988 ();
 FILLCELL_X32 FILLER_123_1009 ();
 FILLCELL_X32 FILLER_123_1041 ();
 FILLCELL_X32 FILLER_123_1073 ();
 FILLCELL_X32 FILLER_123_1105 ();
 FILLCELL_X32 FILLER_123_1137 ();
 FILLCELL_X32 FILLER_123_1169 ();
 FILLCELL_X8 FILLER_123_1201 ();
 FILLCELL_X32 FILLER_124_1 ();
 FILLCELL_X32 FILLER_124_33 ();
 FILLCELL_X32 FILLER_124_65 ();
 FILLCELL_X32 FILLER_124_97 ();
 FILLCELL_X4 FILLER_124_129 ();
 FILLCELL_X8 FILLER_124_143 ();
 FILLCELL_X4 FILLER_124_151 ();
 FILLCELL_X1 FILLER_124_155 ();
 FILLCELL_X2 FILLER_124_163 ();
 FILLCELL_X2 FILLER_124_192 ();
 FILLCELL_X1 FILLER_124_194 ();
 FILLCELL_X16 FILLER_124_197 ();
 FILLCELL_X8 FILLER_124_213 ();
 FILLCELL_X2 FILLER_124_221 ();
 FILLCELL_X1 FILLER_124_223 ();
 FILLCELL_X32 FILLER_124_244 ();
 FILLCELL_X8 FILLER_124_276 ();
 FILLCELL_X4 FILLER_124_284 ();
 FILLCELL_X2 FILLER_124_288 ();
 FILLCELL_X1 FILLER_124_322 ();
 FILLCELL_X8 FILLER_124_340 ();
 FILLCELL_X4 FILLER_124_351 ();
 FILLCELL_X2 FILLER_124_355 ();
 FILLCELL_X1 FILLER_124_362 ();
 FILLCELL_X2 FILLER_124_385 ();
 FILLCELL_X4 FILLER_124_391 ();
 FILLCELL_X2 FILLER_124_395 ();
 FILLCELL_X1 FILLER_124_397 ();
 FILLCELL_X2 FILLER_124_417 ();
 FILLCELL_X1 FILLER_124_419 ();
 FILLCELL_X2 FILLER_124_446 ();
 FILLCELL_X1 FILLER_124_448 ();
 FILLCELL_X16 FILLER_124_463 ();
 FILLCELL_X8 FILLER_124_479 ();
 FILLCELL_X4 FILLER_124_487 ();
 FILLCELL_X2 FILLER_124_532 ();
 FILLCELL_X2 FILLER_124_541 ();
 FILLCELL_X2 FILLER_124_559 ();
 FILLCELL_X16 FILLER_124_567 ();
 FILLCELL_X8 FILLER_124_583 ();
 FILLCELL_X2 FILLER_124_591 ();
 FILLCELL_X1 FILLER_124_593 ();
 FILLCELL_X8 FILLER_124_616 ();
 FILLCELL_X2 FILLER_124_628 ();
 FILLCELL_X1 FILLER_124_630 ();
 FILLCELL_X16 FILLER_124_632 ();
 FILLCELL_X8 FILLER_124_648 ();
 FILLCELL_X4 FILLER_124_656 ();
 FILLCELL_X1 FILLER_124_660 ();
 FILLCELL_X4 FILLER_124_664 ();
 FILLCELL_X2 FILLER_124_668 ();
 FILLCELL_X4 FILLER_124_707 ();
 FILLCELL_X1 FILLER_124_711 ();
 FILLCELL_X16 FILLER_124_734 ();
 FILLCELL_X1 FILLER_124_750 ();
 FILLCELL_X1 FILLER_124_759 ();
 FILLCELL_X2 FILLER_124_772 ();
 FILLCELL_X1 FILLER_124_774 ();
 FILLCELL_X2 FILLER_124_800 ();
 FILLCELL_X8 FILLER_124_807 ();
 FILLCELL_X4 FILLER_124_815 ();
 FILLCELL_X2 FILLER_124_819 ();
 FILLCELL_X2 FILLER_124_845 ();
 FILLCELL_X4 FILLER_124_875 ();
 FILLCELL_X2 FILLER_124_879 ();
 FILLCELL_X1 FILLER_124_901 ();
 FILLCELL_X2 FILLER_124_905 ();
 FILLCELL_X16 FILLER_124_953 ();
 FILLCELL_X4 FILLER_124_969 ();
 FILLCELL_X8 FILLER_124_982 ();
 FILLCELL_X1 FILLER_124_990 ();
 FILLCELL_X8 FILLER_124_1000 ();
 FILLCELL_X2 FILLER_124_1008 ();
 FILLCELL_X1 FILLER_124_1010 ();
 FILLCELL_X16 FILLER_124_1030 ();
 FILLCELL_X2 FILLER_124_1046 ();
 FILLCELL_X1 FILLER_124_1048 ();
 FILLCELL_X32 FILLER_124_1066 ();
 FILLCELL_X32 FILLER_124_1098 ();
 FILLCELL_X32 FILLER_124_1130 ();
 FILLCELL_X32 FILLER_124_1162 ();
 FILLCELL_X8 FILLER_124_1194 ();
 FILLCELL_X4 FILLER_124_1202 ();
 FILLCELL_X2 FILLER_124_1206 ();
 FILLCELL_X1 FILLER_124_1208 ();
 FILLCELL_X32 FILLER_125_1 ();
 FILLCELL_X32 FILLER_125_33 ();
 FILLCELL_X32 FILLER_125_65 ();
 FILLCELL_X32 FILLER_125_97 ();
 FILLCELL_X32 FILLER_125_129 ();
 FILLCELL_X32 FILLER_125_161 ();
 FILLCELL_X1 FILLER_125_193 ();
 FILLCELL_X32 FILLER_125_219 ();
 FILLCELL_X16 FILLER_125_251 ();
 FILLCELL_X8 FILLER_125_267 ();
 FILLCELL_X4 FILLER_125_275 ();
 FILLCELL_X2 FILLER_125_279 ();
 FILLCELL_X8 FILLER_125_327 ();
 FILLCELL_X2 FILLER_125_335 ();
 FILLCELL_X1 FILLER_125_337 ();
 FILLCELL_X1 FILLER_125_358 ();
 FILLCELL_X1 FILLER_125_366 ();
 FILLCELL_X2 FILLER_125_381 ();
 FILLCELL_X1 FILLER_125_383 ();
 FILLCELL_X2 FILLER_125_388 ();
 FILLCELL_X1 FILLER_125_390 ();
 FILLCELL_X4 FILLER_125_403 ();
 FILLCELL_X1 FILLER_125_407 ();
 FILLCELL_X4 FILLER_125_428 ();
 FILLCELL_X1 FILLER_125_432 ();
 FILLCELL_X2 FILLER_125_436 ();
 FILLCELL_X1 FILLER_125_438 ();
 FILLCELL_X4 FILLER_125_444 ();
 FILLCELL_X1 FILLER_125_448 ();
 FILLCELL_X4 FILLER_125_458 ();
 FILLCELL_X1 FILLER_125_462 ();
 FILLCELL_X32 FILLER_125_470 ();
 FILLCELL_X8 FILLER_125_502 ();
 FILLCELL_X8 FILLER_125_532 ();
 FILLCELL_X8 FILLER_125_547 ();
 FILLCELL_X4 FILLER_125_555 ();
 FILLCELL_X2 FILLER_125_559 ();
 FILLCELL_X8 FILLER_125_571 ();
 FILLCELL_X2 FILLER_125_579 ();
 FILLCELL_X4 FILLER_125_583 ();
 FILLCELL_X2 FILLER_125_587 ();
 FILLCELL_X1 FILLER_125_589 ();
 FILLCELL_X4 FILLER_125_602 ();
 FILLCELL_X2 FILLER_125_606 ();
 FILLCELL_X8 FILLER_125_615 ();
 FILLCELL_X1 FILLER_125_623 ();
 FILLCELL_X8 FILLER_125_680 ();
 FILLCELL_X2 FILLER_125_688 ();
 FILLCELL_X1 FILLER_125_690 ();
 FILLCELL_X2 FILLER_125_716 ();
 FILLCELL_X1 FILLER_125_718 ();
 FILLCELL_X16 FILLER_125_729 ();
 FILLCELL_X8 FILLER_125_745 ();
 FILLCELL_X4 FILLER_125_753 ();
 FILLCELL_X1 FILLER_125_761 ();
 FILLCELL_X1 FILLER_125_796 ();
 FILLCELL_X2 FILLER_125_814 ();
 FILLCELL_X2 FILLER_125_831 ();
 FILLCELL_X1 FILLER_125_861 ();
 FILLCELL_X1 FILLER_125_880 ();
 FILLCELL_X8 FILLER_125_885 ();
 FILLCELL_X4 FILLER_125_901 ();
 FILLCELL_X2 FILLER_125_905 ();
 FILLCELL_X1 FILLER_125_914 ();
 FILLCELL_X1 FILLER_125_919 ();
 FILLCELL_X16 FILLER_125_950 ();
 FILLCELL_X4 FILLER_125_966 ();
 FILLCELL_X8 FILLER_125_980 ();
 FILLCELL_X1 FILLER_125_988 ();
 FILLCELL_X32 FILLER_125_999 ();
 FILLCELL_X2 FILLER_125_1031 ();
 FILLCELL_X1 FILLER_125_1033 ();
 FILLCELL_X32 FILLER_125_1053 ();
 FILLCELL_X32 FILLER_125_1085 ();
 FILLCELL_X32 FILLER_125_1117 ();
 FILLCELL_X32 FILLER_125_1149 ();
 FILLCELL_X16 FILLER_125_1181 ();
 FILLCELL_X8 FILLER_125_1197 ();
 FILLCELL_X4 FILLER_125_1205 ();
 FILLCELL_X32 FILLER_126_1 ();
 FILLCELL_X32 FILLER_126_33 ();
 FILLCELL_X32 FILLER_126_65 ();
 FILLCELL_X32 FILLER_126_97 ();
 FILLCELL_X32 FILLER_126_129 ();
 FILLCELL_X32 FILLER_126_161 ();
 FILLCELL_X32 FILLER_126_193 ();
 FILLCELL_X32 FILLER_126_225 ();
 FILLCELL_X16 FILLER_126_257 ();
 FILLCELL_X4 FILLER_126_273 ();
 FILLCELL_X1 FILLER_126_277 ();
 FILLCELL_X2 FILLER_126_330 ();
 FILLCELL_X1 FILLER_126_332 ();
 FILLCELL_X8 FILLER_126_340 ();
 FILLCELL_X2 FILLER_126_361 ();
 FILLCELL_X2 FILLER_126_386 ();
 FILLCELL_X1 FILLER_126_388 ();
 FILLCELL_X1 FILLER_126_405 ();
 FILLCELL_X1 FILLER_126_410 ();
 FILLCELL_X2 FILLER_126_431 ();
 FILLCELL_X1 FILLER_126_433 ();
 FILLCELL_X4 FILLER_126_441 ();
 FILLCELL_X32 FILLER_126_453 ();
 FILLCELL_X8 FILLER_126_485 ();
 FILLCELL_X2 FILLER_126_522 ();
 FILLCELL_X1 FILLER_126_524 ();
 FILLCELL_X2 FILLER_126_552 ();
 FILLCELL_X2 FILLER_126_573 ();
 FILLCELL_X4 FILLER_126_581 ();
 FILLCELL_X1 FILLER_126_585 ();
 FILLCELL_X1 FILLER_126_609 ();
 FILLCELL_X4 FILLER_126_627 ();
 FILLCELL_X8 FILLER_126_645 ();
 FILLCELL_X2 FILLER_126_653 ();
 FILLCELL_X2 FILLER_126_672 ();
 FILLCELL_X1 FILLER_126_674 ();
 FILLCELL_X8 FILLER_126_681 ();
 FILLCELL_X2 FILLER_126_689 ();
 FILLCELL_X4 FILLER_126_714 ();
 FILLCELL_X1 FILLER_126_735 ();
 FILLCELL_X8 FILLER_126_741 ();
 FILLCELL_X1 FILLER_126_749 ();
 FILLCELL_X1 FILLER_126_764 ();
 FILLCELL_X2 FILLER_126_772 ();
 FILLCELL_X1 FILLER_126_791 ();
 FILLCELL_X1 FILLER_126_828 ();
 FILLCELL_X4 FILLER_126_844 ();
 FILLCELL_X1 FILLER_126_848 ();
 FILLCELL_X2 FILLER_126_876 ();
 FILLCELL_X2 FILLER_126_885 ();
 FILLCELL_X1 FILLER_126_887 ();
 FILLCELL_X8 FILLER_126_896 ();
 FILLCELL_X4 FILLER_126_904 ();
 FILLCELL_X1 FILLER_126_908 ();
 FILLCELL_X16 FILLER_126_953 ();
 FILLCELL_X8 FILLER_126_969 ();
 FILLCELL_X16 FILLER_126_990 ();
 FILLCELL_X4 FILLER_126_1006 ();
 FILLCELL_X2 FILLER_126_1010 ();
 FILLCELL_X1 FILLER_126_1012 ();
 FILLCELL_X2 FILLER_126_1020 ();
 FILLCELL_X4 FILLER_126_1029 ();
 FILLCELL_X2 FILLER_126_1033 ();
 FILLCELL_X32 FILLER_126_1063 ();
 FILLCELL_X32 FILLER_126_1095 ();
 FILLCELL_X32 FILLER_126_1127 ();
 FILLCELL_X32 FILLER_126_1159 ();
 FILLCELL_X16 FILLER_126_1191 ();
 FILLCELL_X2 FILLER_126_1207 ();
 FILLCELL_X32 FILLER_127_1 ();
 FILLCELL_X32 FILLER_127_33 ();
 FILLCELL_X32 FILLER_127_65 ();
 FILLCELL_X32 FILLER_127_97 ();
 FILLCELL_X32 FILLER_127_129 ();
 FILLCELL_X32 FILLER_127_161 ();
 FILLCELL_X32 FILLER_127_193 ();
 FILLCELL_X32 FILLER_127_225 ();
 FILLCELL_X1 FILLER_127_257 ();
 FILLCELL_X2 FILLER_127_334 ();
 FILLCELL_X2 FILLER_127_347 ();
 FILLCELL_X16 FILLER_127_401 ();
 FILLCELL_X2 FILLER_127_417 ();
 FILLCELL_X1 FILLER_127_419 ();
 FILLCELL_X2 FILLER_127_436 ();
 FILLCELL_X1 FILLER_127_446 ();
 FILLCELL_X4 FILLER_127_451 ();
 FILLCELL_X16 FILLER_127_460 ();
 FILLCELL_X2 FILLER_127_476 ();
 FILLCELL_X4 FILLER_127_495 ();
 FILLCELL_X2 FILLER_127_499 ();
 FILLCELL_X1 FILLER_127_501 ();
 FILLCELL_X2 FILLER_127_519 ();
 FILLCELL_X1 FILLER_127_521 ();
 FILLCELL_X1 FILLER_127_532 ();
 FILLCELL_X1 FILLER_127_580 ();
 FILLCELL_X1 FILLER_127_606 ();
 FILLCELL_X4 FILLER_127_634 ();
 FILLCELL_X1 FILLER_127_669 ();
 FILLCELL_X1 FILLER_127_677 ();
 FILLCELL_X1 FILLER_127_695 ();
 FILLCELL_X2 FILLER_127_702 ();
 FILLCELL_X2 FILLER_127_710 ();
 FILLCELL_X2 FILLER_127_718 ();
 FILLCELL_X16 FILLER_127_727 ();
 FILLCELL_X8 FILLER_127_743 ();
 FILLCELL_X4 FILLER_127_751 ();
 FILLCELL_X2 FILLER_127_755 ();
 FILLCELL_X1 FILLER_127_757 ();
 FILLCELL_X2 FILLER_127_763 ();
 FILLCELL_X2 FILLER_127_770 ();
 FILLCELL_X1 FILLER_127_772 ();
 FILLCELL_X2 FILLER_127_777 ();
 FILLCELL_X1 FILLER_127_795 ();
 FILLCELL_X1 FILLER_127_807 ();
 FILLCELL_X4 FILLER_127_815 ();
 FILLCELL_X2 FILLER_127_819 ();
 FILLCELL_X1 FILLER_127_821 ();
 FILLCELL_X2 FILLER_127_827 ();
 FILLCELL_X1 FILLER_127_829 ();
 FILLCELL_X1 FILLER_127_839 ();
 FILLCELL_X1 FILLER_127_862 ();
 FILLCELL_X4 FILLER_127_867 ();
 FILLCELL_X2 FILLER_127_871 ();
 FILLCELL_X4 FILLER_127_876 ();
 FILLCELL_X16 FILLER_127_884 ();
 FILLCELL_X2 FILLER_127_900 ();
 FILLCELL_X1 FILLER_127_902 ();
 FILLCELL_X4 FILLER_127_926 ();
 FILLCELL_X4 FILLER_127_940 ();
 FILLCELL_X16 FILLER_127_951 ();
 FILLCELL_X8 FILLER_127_967 ();
 FILLCELL_X4 FILLER_127_975 ();
 FILLCELL_X2 FILLER_127_995 ();
 FILLCELL_X2 FILLER_127_1004 ();
 FILLCELL_X2 FILLER_127_1011 ();
 FILLCELL_X1 FILLER_127_1013 ();
 FILLCELL_X4 FILLER_127_1021 ();
 FILLCELL_X2 FILLER_127_1030 ();
 FILLCELL_X32 FILLER_127_1082 ();
 FILLCELL_X32 FILLER_127_1114 ();
 FILLCELL_X32 FILLER_127_1146 ();
 FILLCELL_X16 FILLER_127_1178 ();
 FILLCELL_X8 FILLER_127_1194 ();
 FILLCELL_X4 FILLER_127_1202 ();
 FILLCELL_X2 FILLER_127_1206 ();
 FILLCELL_X1 FILLER_127_1208 ();
 FILLCELL_X32 FILLER_128_1 ();
 FILLCELL_X32 FILLER_128_33 ();
 FILLCELL_X32 FILLER_128_65 ();
 FILLCELL_X32 FILLER_128_97 ();
 FILLCELL_X32 FILLER_128_129 ();
 FILLCELL_X32 FILLER_128_161 ();
 FILLCELL_X32 FILLER_128_193 ();
 FILLCELL_X32 FILLER_128_225 ();
 FILLCELL_X8 FILLER_128_257 ();
 FILLCELL_X2 FILLER_128_265 ();
 FILLCELL_X2 FILLER_128_280 ();
 FILLCELL_X2 FILLER_128_312 ();
 FILLCELL_X1 FILLER_128_314 ();
 FILLCELL_X1 FILLER_128_320 ();
 FILLCELL_X1 FILLER_128_328 ();
 FILLCELL_X2 FILLER_128_335 ();
 FILLCELL_X1 FILLER_128_370 ();
 FILLCELL_X2 FILLER_128_385 ();
 FILLCELL_X1 FILLER_128_387 ();
 FILLCELL_X2 FILLER_128_438 ();
 FILLCELL_X8 FILLER_128_463 ();
 FILLCELL_X4 FILLER_128_471 ();
 FILLCELL_X2 FILLER_128_475 ();
 FILLCELL_X16 FILLER_128_480 ();
 FILLCELL_X1 FILLER_128_496 ();
 FILLCELL_X1 FILLER_128_532 ();
 FILLCELL_X2 FILLER_128_539 ();
 FILLCELL_X1 FILLER_128_541 ();
 FILLCELL_X8 FILLER_128_546 ();
 FILLCELL_X1 FILLER_128_554 ();
 FILLCELL_X2 FILLER_128_583 ();
 FILLCELL_X2 FILLER_128_591 ();
 FILLCELL_X4 FILLER_128_624 ();
 FILLCELL_X2 FILLER_128_628 ();
 FILLCELL_X1 FILLER_128_630 ();
 FILLCELL_X2 FILLER_128_632 ();
 FILLCELL_X4 FILLER_128_641 ();
 FILLCELL_X1 FILLER_128_645 ();
 FILLCELL_X4 FILLER_128_654 ();
 FILLCELL_X16 FILLER_128_666 ();
 FILLCELL_X4 FILLER_128_682 ();
 FILLCELL_X4 FILLER_128_698 ();
 FILLCELL_X2 FILLER_128_702 ();
 FILLCELL_X2 FILLER_128_720 ();
 FILLCELL_X16 FILLER_128_744 ();
 FILLCELL_X8 FILLER_128_760 ();
 FILLCELL_X2 FILLER_128_768 ();
 FILLCELL_X4 FILLER_128_774 ();
 FILLCELL_X2 FILLER_128_778 ();
 FILLCELL_X1 FILLER_128_780 ();
 FILLCELL_X2 FILLER_128_809 ();
 FILLCELL_X1 FILLER_128_811 ();
 FILLCELL_X1 FILLER_128_824 ();
 FILLCELL_X2 FILLER_128_839 ();
 FILLCELL_X1 FILLER_128_841 ();
 FILLCELL_X4 FILLER_128_846 ();
 FILLCELL_X2 FILLER_128_857 ();
 FILLCELL_X1 FILLER_128_864 ();
 FILLCELL_X1 FILLER_128_876 ();
 FILLCELL_X2 FILLER_128_901 ();
 FILLCELL_X2 FILLER_128_929 ();
 FILLCELL_X16 FILLER_128_944 ();
 FILLCELL_X8 FILLER_128_960 ();
 FILLCELL_X4 FILLER_128_968 ();
 FILLCELL_X2 FILLER_128_972 ();
 FILLCELL_X4 FILLER_128_991 ();
 FILLCELL_X1 FILLER_128_1031 ();
 FILLCELL_X1 FILLER_128_1041 ();
 FILLCELL_X2 FILLER_128_1057 ();
 FILLCELL_X32 FILLER_128_1086 ();
 FILLCELL_X32 FILLER_128_1118 ();
 FILLCELL_X32 FILLER_128_1150 ();
 FILLCELL_X16 FILLER_128_1182 ();
 FILLCELL_X8 FILLER_128_1198 ();
 FILLCELL_X2 FILLER_128_1206 ();
 FILLCELL_X1 FILLER_128_1208 ();
 FILLCELL_X32 FILLER_129_1 ();
 FILLCELL_X32 FILLER_129_33 ();
 FILLCELL_X32 FILLER_129_65 ();
 FILLCELL_X32 FILLER_129_97 ();
 FILLCELL_X32 FILLER_129_129 ();
 FILLCELL_X32 FILLER_129_161 ();
 FILLCELL_X32 FILLER_129_193 ();
 FILLCELL_X32 FILLER_129_225 ();
 FILLCELL_X32 FILLER_129_257 ();
 FILLCELL_X2 FILLER_129_302 ();
 FILLCELL_X2 FILLER_129_389 ();
 FILLCELL_X1 FILLER_129_391 ();
 FILLCELL_X1 FILLER_129_401 ();
 FILLCELL_X2 FILLER_129_413 ();
 FILLCELL_X1 FILLER_129_415 ();
 FILLCELL_X1 FILLER_129_432 ();
 FILLCELL_X8 FILLER_129_459 ();
 FILLCELL_X1 FILLER_129_467 ();
 FILLCELL_X8 FILLER_129_475 ();
 FILLCELL_X1 FILLER_129_483 ();
 FILLCELL_X16 FILLER_129_501 ();
 FILLCELL_X4 FILLER_129_530 ();
 FILLCELL_X2 FILLER_129_534 ();
 FILLCELL_X2 FILLER_129_542 ();
 FILLCELL_X2 FILLER_129_551 ();
 FILLCELL_X1 FILLER_129_553 ();
 FILLCELL_X1 FILLER_129_572 ();
 FILLCELL_X2 FILLER_129_585 ();
 FILLCELL_X8 FILLER_129_594 ();
 FILLCELL_X2 FILLER_129_602 ();
 FILLCELL_X1 FILLER_129_604 ();
 FILLCELL_X1 FILLER_129_624 ();
 FILLCELL_X2 FILLER_129_653 ();
 FILLCELL_X1 FILLER_129_655 ();
 FILLCELL_X16 FILLER_129_660 ();
 FILLCELL_X8 FILLER_129_676 ();
 FILLCELL_X1 FILLER_129_705 ();
 FILLCELL_X1 FILLER_129_715 ();
 FILLCELL_X16 FILLER_129_723 ();
 FILLCELL_X4 FILLER_129_739 ();
 FILLCELL_X2 FILLER_129_743 ();
 FILLCELL_X16 FILLER_129_752 ();
 FILLCELL_X2 FILLER_129_768 ();
 FILLCELL_X8 FILLER_129_783 ();
 FILLCELL_X1 FILLER_129_791 ();
 FILLCELL_X1 FILLER_129_798 ();
 FILLCELL_X2 FILLER_129_815 ();
 FILLCELL_X1 FILLER_129_817 ();
 FILLCELL_X2 FILLER_129_827 ();
 FILLCELL_X1 FILLER_129_829 ();
 FILLCELL_X4 FILLER_129_837 ();
 FILLCELL_X1 FILLER_129_841 ();
 FILLCELL_X2 FILLER_129_852 ();
 FILLCELL_X4 FILLER_129_857 ();
 FILLCELL_X2 FILLER_129_887 ();
 FILLCELL_X4 FILLER_129_899 ();
 FILLCELL_X32 FILLER_129_910 ();
 FILLCELL_X16 FILLER_129_942 ();
 FILLCELL_X4 FILLER_129_958 ();
 FILLCELL_X2 FILLER_129_978 ();
 FILLCELL_X4 FILLER_129_1031 ();
 FILLCELL_X1 FILLER_129_1035 ();
 FILLCELL_X1 FILLER_129_1050 ();
 FILLCELL_X1 FILLER_129_1055 ();
 FILLCELL_X2 FILLER_129_1084 ();
 FILLCELL_X32 FILLER_129_1093 ();
 FILLCELL_X32 FILLER_129_1125 ();
 FILLCELL_X32 FILLER_129_1157 ();
 FILLCELL_X16 FILLER_129_1189 ();
 FILLCELL_X4 FILLER_129_1205 ();
 FILLCELL_X32 FILLER_130_1 ();
 FILLCELL_X32 FILLER_130_33 ();
 FILLCELL_X32 FILLER_130_65 ();
 FILLCELL_X32 FILLER_130_97 ();
 FILLCELL_X32 FILLER_130_129 ();
 FILLCELL_X32 FILLER_130_161 ();
 FILLCELL_X32 FILLER_130_193 ();
 FILLCELL_X32 FILLER_130_225 ();
 FILLCELL_X16 FILLER_130_257 ();
 FILLCELL_X4 FILLER_130_286 ();
 FILLCELL_X2 FILLER_130_339 ();
 FILLCELL_X8 FILLER_130_349 ();
 FILLCELL_X4 FILLER_130_357 ();
 FILLCELL_X2 FILLER_130_361 ();
 FILLCELL_X1 FILLER_130_363 ();
 FILLCELL_X1 FILLER_130_393 ();
 FILLCELL_X4 FILLER_130_411 ();
 FILLCELL_X1 FILLER_130_415 ();
 FILLCELL_X2 FILLER_130_430 ();
 FILLCELL_X1 FILLER_130_435 ();
 FILLCELL_X2 FILLER_130_440 ();
 FILLCELL_X1 FILLER_130_442 ();
 FILLCELL_X32 FILLER_130_448 ();
 FILLCELL_X2 FILLER_130_480 ();
 FILLCELL_X1 FILLER_130_482 ();
 FILLCELL_X8 FILLER_130_500 ();
 FILLCELL_X2 FILLER_130_508 ();
 FILLCELL_X1 FILLER_130_510 ();
 FILLCELL_X8 FILLER_130_527 ();
 FILLCELL_X2 FILLER_130_542 ();
 FILLCELL_X1 FILLER_130_544 ();
 FILLCELL_X4 FILLER_130_562 ();
 FILLCELL_X2 FILLER_130_566 ();
 FILLCELL_X4 FILLER_130_575 ();
 FILLCELL_X2 FILLER_130_579 ();
 FILLCELL_X1 FILLER_130_581 ();
 FILLCELL_X2 FILLER_130_592 ();
 FILLCELL_X1 FILLER_130_607 ();
 FILLCELL_X1 FILLER_130_621 ();
 FILLCELL_X32 FILLER_130_706 ();
 FILLCELL_X2 FILLER_130_738 ();
 FILLCELL_X1 FILLER_130_740 ();
 FILLCELL_X32 FILLER_130_750 ();
 FILLCELL_X8 FILLER_130_782 ();
 FILLCELL_X4 FILLER_130_790 ();
 FILLCELL_X2 FILLER_130_794 ();
 FILLCELL_X1 FILLER_130_803 ();
 FILLCELL_X4 FILLER_130_817 ();
 FILLCELL_X2 FILLER_130_821 ();
 FILLCELL_X4 FILLER_130_833 ();
 FILLCELL_X8 FILLER_130_854 ();
 FILLCELL_X2 FILLER_130_862 ();
 FILLCELL_X2 FILLER_130_876 ();
 FILLCELL_X1 FILLER_130_878 ();
 FILLCELL_X32 FILLER_130_898 ();
 FILLCELL_X4 FILLER_130_930 ();
 FILLCELL_X1 FILLER_130_934 ();
 FILLCELL_X2 FILLER_130_940 ();
 FILLCELL_X2 FILLER_130_956 ();
 FILLCELL_X1 FILLER_130_958 ();
 FILLCELL_X2 FILLER_130_1028 ();
 FILLCELL_X1 FILLER_130_1030 ();
 FILLCELL_X1 FILLER_130_1038 ();
 FILLCELL_X4 FILLER_130_1045 ();
 FILLCELL_X2 FILLER_130_1049 ();
 FILLCELL_X2 FILLER_130_1076 ();
 FILLCELL_X32 FILLER_130_1088 ();
 FILLCELL_X32 FILLER_130_1120 ();
 FILLCELL_X32 FILLER_130_1152 ();
 FILLCELL_X16 FILLER_130_1184 ();
 FILLCELL_X8 FILLER_130_1200 ();
 FILLCELL_X1 FILLER_130_1208 ();
 FILLCELL_X32 FILLER_131_1 ();
 FILLCELL_X32 FILLER_131_33 ();
 FILLCELL_X32 FILLER_131_65 ();
 FILLCELL_X32 FILLER_131_97 ();
 FILLCELL_X32 FILLER_131_129 ();
 FILLCELL_X32 FILLER_131_161 ();
 FILLCELL_X32 FILLER_131_193 ();
 FILLCELL_X32 FILLER_131_225 ();
 FILLCELL_X8 FILLER_131_257 ();
 FILLCELL_X4 FILLER_131_265 ();
 FILLCELL_X2 FILLER_131_269 ();
 FILLCELL_X4 FILLER_131_298 ();
 FILLCELL_X1 FILLER_131_302 ();
 FILLCELL_X4 FILLER_131_317 ();
 FILLCELL_X8 FILLER_131_334 ();
 FILLCELL_X4 FILLER_131_342 ();
 FILLCELL_X4 FILLER_131_359 ();
 FILLCELL_X2 FILLER_131_363 ();
 FILLCELL_X1 FILLER_131_365 ();
 FILLCELL_X2 FILLER_131_373 ();
 FILLCELL_X1 FILLER_131_375 ();
 FILLCELL_X8 FILLER_131_403 ();
 FILLCELL_X4 FILLER_131_411 ();
 FILLCELL_X2 FILLER_131_415 ();
 FILLCELL_X1 FILLER_131_417 ();
 FILLCELL_X2 FILLER_131_422 ();
 FILLCELL_X1 FILLER_131_424 ();
 FILLCELL_X8 FILLER_131_444 ();
 FILLCELL_X4 FILLER_131_452 ();
 FILLCELL_X1 FILLER_131_456 ();
 FILLCELL_X4 FILLER_131_474 ();
 FILLCELL_X32 FILLER_131_506 ();
 FILLCELL_X16 FILLER_131_538 ();
 FILLCELL_X2 FILLER_131_554 ();
 FILLCELL_X1 FILLER_131_556 ();
 FILLCELL_X2 FILLER_131_570 ();
 FILLCELL_X2 FILLER_131_589 ();
 FILLCELL_X1 FILLER_131_591 ();
 FILLCELL_X2 FILLER_131_637 ();
 FILLCELL_X2 FILLER_131_658 ();
 FILLCELL_X16 FILLER_131_667 ();
 FILLCELL_X8 FILLER_131_683 ();
 FILLCELL_X4 FILLER_131_691 ();
 FILLCELL_X2 FILLER_131_695 ();
 FILLCELL_X1 FILLER_131_697 ();
 FILLCELL_X2 FILLER_131_715 ();
 FILLCELL_X2 FILLER_131_726 ();
 FILLCELL_X1 FILLER_131_728 ();
 FILLCELL_X16 FILLER_131_747 ();
 FILLCELL_X4 FILLER_131_763 ();
 FILLCELL_X2 FILLER_131_767 ();
 FILLCELL_X1 FILLER_131_769 ();
 FILLCELL_X2 FILLER_131_786 ();
 FILLCELL_X32 FILLER_131_795 ();
 FILLCELL_X32 FILLER_131_827 ();
 FILLCELL_X8 FILLER_131_859 ();
 FILLCELL_X4 FILLER_131_867 ();
 FILLCELL_X2 FILLER_131_871 ();
 FILLCELL_X4 FILLER_131_883 ();
 FILLCELL_X1 FILLER_131_887 ();
 FILLCELL_X16 FILLER_131_907 ();
 FILLCELL_X8 FILLER_131_923 ();
 FILLCELL_X2 FILLER_131_931 ();
 FILLCELL_X8 FILLER_131_954 ();
 FILLCELL_X4 FILLER_131_962 ();
 FILLCELL_X2 FILLER_131_966 ();
 FILLCELL_X1 FILLER_131_968 ();
 FILLCELL_X2 FILLER_131_994 ();
 FILLCELL_X1 FILLER_131_1008 ();
 FILLCELL_X1 FILLER_131_1023 ();
 FILLCELL_X2 FILLER_131_1035 ();
 FILLCELL_X2 FILLER_131_1055 ();
 FILLCELL_X1 FILLER_131_1057 ();
 FILLCELL_X4 FILLER_131_1061 ();
 FILLCELL_X2 FILLER_131_1065 ();
 FILLCELL_X1 FILLER_131_1067 ();
 FILLCELL_X2 FILLER_131_1071 ();
 FILLCELL_X1 FILLER_131_1073 ();
 FILLCELL_X1 FILLER_131_1082 ();
 FILLCELL_X2 FILLER_131_1087 ();
 FILLCELL_X1 FILLER_131_1089 ();
 FILLCELL_X2 FILLER_131_1094 ();
 FILLCELL_X1 FILLER_131_1096 ();
 FILLCELL_X32 FILLER_131_1118 ();
 FILLCELL_X32 FILLER_131_1150 ();
 FILLCELL_X16 FILLER_131_1182 ();
 FILLCELL_X8 FILLER_131_1198 ();
 FILLCELL_X2 FILLER_131_1206 ();
 FILLCELL_X1 FILLER_131_1208 ();
 FILLCELL_X32 FILLER_132_1 ();
 FILLCELL_X32 FILLER_132_33 ();
 FILLCELL_X32 FILLER_132_65 ();
 FILLCELL_X32 FILLER_132_97 ();
 FILLCELL_X32 FILLER_132_129 ();
 FILLCELL_X32 FILLER_132_161 ();
 FILLCELL_X32 FILLER_132_193 ();
 FILLCELL_X16 FILLER_132_225 ();
 FILLCELL_X8 FILLER_132_241 ();
 FILLCELL_X4 FILLER_132_249 ();
 FILLCELL_X2 FILLER_132_253 ();
 FILLCELL_X2 FILLER_132_278 ();
 FILLCELL_X1 FILLER_132_280 ();
 FILLCELL_X4 FILLER_132_301 ();
 FILLCELL_X4 FILLER_132_318 ();
 FILLCELL_X2 FILLER_132_322 ();
 FILLCELL_X1 FILLER_132_324 ();
 FILLCELL_X2 FILLER_132_338 ();
 FILLCELL_X1 FILLER_132_353 ();
 FILLCELL_X16 FILLER_132_361 ();
 FILLCELL_X2 FILLER_132_377 ();
 FILLCELL_X1 FILLER_132_379 ();
 FILLCELL_X1 FILLER_132_384 ();
 FILLCELL_X16 FILLER_132_396 ();
 FILLCELL_X4 FILLER_132_412 ();
 FILLCELL_X2 FILLER_132_416 ();
 FILLCELL_X16 FILLER_132_425 ();
 FILLCELL_X4 FILLER_132_441 ();
 FILLCELL_X1 FILLER_132_445 ();
 FILLCELL_X16 FILLER_132_468 ();
 FILLCELL_X2 FILLER_132_484 ();
 FILLCELL_X1 FILLER_132_486 ();
 FILLCELL_X16 FILLER_132_506 ();
 FILLCELL_X1 FILLER_132_522 ();
 FILLCELL_X1 FILLER_132_537 ();
 FILLCELL_X8 FILLER_132_547 ();
 FILLCELL_X4 FILLER_132_555 ();
 FILLCELL_X2 FILLER_132_559 ();
 FILLCELL_X1 FILLER_132_561 ();
 FILLCELL_X16 FILLER_132_604 ();
 FILLCELL_X2 FILLER_132_620 ();
 FILLCELL_X1 FILLER_132_622 ();
 FILLCELL_X4 FILLER_132_627 ();
 FILLCELL_X8 FILLER_132_632 ();
 FILLCELL_X2 FILLER_132_640 ();
 FILLCELL_X1 FILLER_132_642 ();
 FILLCELL_X1 FILLER_132_645 ();
 FILLCELL_X1 FILLER_132_649 ();
 FILLCELL_X4 FILLER_132_667 ();
 FILLCELL_X8 FILLER_132_677 ();
 FILLCELL_X4 FILLER_132_699 ();
 FILLCELL_X2 FILLER_132_703 ();
 FILLCELL_X1 FILLER_132_705 ();
 FILLCELL_X2 FILLER_132_736 ();
 FILLCELL_X1 FILLER_132_738 ();
 FILLCELL_X8 FILLER_132_760 ();
 FILLCELL_X4 FILLER_132_768 ();
 FILLCELL_X32 FILLER_132_789 ();
 FILLCELL_X8 FILLER_132_821 ();
 FILLCELL_X4 FILLER_132_829 ();
 FILLCELL_X2 FILLER_132_833 ();
 FILLCELL_X8 FILLER_132_857 ();
 FILLCELL_X4 FILLER_132_865 ();
 FILLCELL_X8 FILLER_132_875 ();
 FILLCELL_X4 FILLER_132_883 ();
 FILLCELL_X1 FILLER_132_887 ();
 FILLCELL_X4 FILLER_132_937 ();
 FILLCELL_X1 FILLER_132_941 ();
 FILLCELL_X4 FILLER_132_963 ();
 FILLCELL_X1 FILLER_132_974 ();
 FILLCELL_X2 FILLER_132_985 ();
 FILLCELL_X1 FILLER_132_1002 ();
 FILLCELL_X1 FILLER_132_1020 ();
 FILLCELL_X2 FILLER_132_1028 ();
 FILLCELL_X4 FILLER_132_1086 ();
 FILLCELL_X2 FILLER_132_1090 ();
 FILLCELL_X1 FILLER_132_1092 ();
 FILLCELL_X8 FILLER_132_1108 ();
 FILLCELL_X32 FILLER_132_1126 ();
 FILLCELL_X32 FILLER_132_1158 ();
 FILLCELL_X16 FILLER_132_1190 ();
 FILLCELL_X2 FILLER_132_1206 ();
 FILLCELL_X1 FILLER_132_1208 ();
 FILLCELL_X32 FILLER_133_1 ();
 FILLCELL_X32 FILLER_133_33 ();
 FILLCELL_X32 FILLER_133_65 ();
 FILLCELL_X32 FILLER_133_97 ();
 FILLCELL_X32 FILLER_133_129 ();
 FILLCELL_X32 FILLER_133_161 ();
 FILLCELL_X32 FILLER_133_193 ();
 FILLCELL_X4 FILLER_133_225 ();
 FILLCELL_X8 FILLER_133_242 ();
 FILLCELL_X1 FILLER_133_250 ();
 FILLCELL_X1 FILLER_133_267 ();
 FILLCELL_X8 FILLER_133_287 ();
 FILLCELL_X4 FILLER_133_295 ();
 FILLCELL_X2 FILLER_133_312 ();
 FILLCELL_X1 FILLER_133_314 ();
 FILLCELL_X2 FILLER_133_348 ();
 FILLCELL_X32 FILLER_133_397 ();
 FILLCELL_X4 FILLER_133_429 ();
 FILLCELL_X2 FILLER_133_433 ();
 FILLCELL_X16 FILLER_133_459 ();
 FILLCELL_X4 FILLER_133_478 ();
 FILLCELL_X2 FILLER_133_482 ();
 FILLCELL_X8 FILLER_133_494 ();
 FILLCELL_X4 FILLER_133_502 ();
 FILLCELL_X4 FILLER_133_513 ();
 FILLCELL_X1 FILLER_133_517 ();
 FILLCELL_X4 FILLER_133_525 ();
 FILLCELL_X4 FILLER_133_532 ();
 FILLCELL_X8 FILLER_133_550 ();
 FILLCELL_X2 FILLER_133_558 ();
 FILLCELL_X1 FILLER_133_560 ();
 FILLCELL_X8 FILLER_133_564 ();
 FILLCELL_X2 FILLER_133_572 ();
 FILLCELL_X1 FILLER_133_580 ();
 FILLCELL_X4 FILLER_133_589 ();
 FILLCELL_X2 FILLER_133_593 ();
 FILLCELL_X32 FILLER_133_604 ();
 FILLCELL_X32 FILLER_133_636 ();
 FILLCELL_X4 FILLER_133_668 ();
 FILLCELL_X16 FILLER_133_689 ();
 FILLCELL_X4 FILLER_133_705 ();
 FILLCELL_X4 FILLER_133_740 ();
 FILLCELL_X2 FILLER_133_744 ();
 FILLCELL_X1 FILLER_133_746 ();
 FILLCELL_X16 FILLER_133_761 ();
 FILLCELL_X4 FILLER_133_777 ();
 FILLCELL_X2 FILLER_133_781 ();
 FILLCELL_X1 FILLER_133_783 ();
 FILLCELL_X4 FILLER_133_806 ();
 FILLCELL_X16 FILLER_133_827 ();
 FILLCELL_X8 FILLER_133_843 ();
 FILLCELL_X2 FILLER_133_851 ();
 FILLCELL_X8 FILLER_133_859 ();
 FILLCELL_X2 FILLER_133_867 ();
 FILLCELL_X1 FILLER_133_869 ();
 FILLCELL_X16 FILLER_133_887 ();
 FILLCELL_X4 FILLER_133_903 ();
 FILLCELL_X2 FILLER_133_907 ();
 FILLCELL_X2 FILLER_133_916 ();
 FILLCELL_X1 FILLER_133_918 ();
 FILLCELL_X1 FILLER_133_922 ();
 FILLCELL_X4 FILLER_133_926 ();
 FILLCELL_X2 FILLER_133_930 ();
 FILLCELL_X2 FILLER_133_950 ();
 FILLCELL_X1 FILLER_133_952 ();
 FILLCELL_X2 FILLER_133_960 ();
 FILLCELL_X1 FILLER_133_979 ();
 FILLCELL_X2 FILLER_133_987 ();
 FILLCELL_X1 FILLER_133_1001 ();
 FILLCELL_X2 FILLER_133_1006 ();
 FILLCELL_X2 FILLER_133_1026 ();
 FILLCELL_X1 FILLER_133_1032 ();
 FILLCELL_X4 FILLER_133_1070 ();
 FILLCELL_X2 FILLER_133_1074 ();
 FILLCELL_X1 FILLER_133_1076 ();
 FILLCELL_X4 FILLER_133_1081 ();
 FILLCELL_X2 FILLER_133_1085 ();
 FILLCELL_X1 FILLER_133_1087 ();
 FILLCELL_X2 FILLER_133_1111 ();
 FILLCELL_X1 FILLER_133_1120 ();
 FILLCELL_X32 FILLER_133_1125 ();
 FILLCELL_X32 FILLER_133_1157 ();
 FILLCELL_X16 FILLER_133_1189 ();
 FILLCELL_X4 FILLER_133_1205 ();
 FILLCELL_X32 FILLER_134_1 ();
 FILLCELL_X32 FILLER_134_33 ();
 FILLCELL_X32 FILLER_134_65 ();
 FILLCELL_X32 FILLER_134_97 ();
 FILLCELL_X32 FILLER_134_129 ();
 FILLCELL_X32 FILLER_134_161 ();
 FILLCELL_X32 FILLER_134_193 ();
 FILLCELL_X1 FILLER_134_225 ();
 FILLCELL_X4 FILLER_134_245 ();
 FILLCELL_X2 FILLER_134_249 ();
 FILLCELL_X2 FILLER_134_258 ();
 FILLCELL_X1 FILLER_134_293 ();
 FILLCELL_X2 FILLER_134_339 ();
 FILLCELL_X8 FILLER_134_388 ();
 FILLCELL_X2 FILLER_134_396 ();
 FILLCELL_X1 FILLER_134_398 ();
 FILLCELL_X8 FILLER_134_446 ();
 FILLCELL_X4 FILLER_134_454 ();
 FILLCELL_X4 FILLER_134_465 ();
 FILLCELL_X2 FILLER_134_488 ();
 FILLCELL_X8 FILLER_134_511 ();
 FILLCELL_X1 FILLER_134_519 ();
 FILLCELL_X8 FILLER_134_548 ();
 FILLCELL_X4 FILLER_134_556 ();
 FILLCELL_X2 FILLER_134_560 ();
 FILLCELL_X4 FILLER_134_568 ();
 FILLCELL_X4 FILLER_134_577 ();
 FILLCELL_X2 FILLER_134_581 ();
 FILLCELL_X1 FILLER_134_583 ();
 FILLCELL_X16 FILLER_134_610 ();
 FILLCELL_X4 FILLER_134_626 ();
 FILLCELL_X1 FILLER_134_630 ();
 FILLCELL_X8 FILLER_134_632 ();
 FILLCELL_X4 FILLER_134_640 ();
 FILLCELL_X1 FILLER_134_644 ();
 FILLCELL_X2 FILLER_134_652 ();
 FILLCELL_X16 FILLER_134_662 ();
 FILLCELL_X8 FILLER_134_678 ();
 FILLCELL_X4 FILLER_134_686 ();
 FILLCELL_X8 FILLER_134_704 ();
 FILLCELL_X16 FILLER_134_729 ();
 FILLCELL_X4 FILLER_134_745 ();
 FILLCELL_X2 FILLER_134_749 ();
 FILLCELL_X4 FILLER_134_768 ();
 FILLCELL_X2 FILLER_134_772 ();
 FILLCELL_X1 FILLER_134_774 ();
 FILLCELL_X2 FILLER_134_780 ();
 FILLCELL_X1 FILLER_134_782 ();
 FILLCELL_X32 FILLER_134_790 ();
 FILLCELL_X2 FILLER_134_822 ();
 FILLCELL_X1 FILLER_134_824 ();
 FILLCELL_X8 FILLER_134_832 ();
 FILLCELL_X2 FILLER_134_840 ();
 FILLCELL_X1 FILLER_134_842 ();
 FILLCELL_X4 FILLER_134_847 ();
 FILLCELL_X2 FILLER_134_851 ();
 FILLCELL_X8 FILLER_134_878 ();
 FILLCELL_X1 FILLER_134_886 ();
 FILLCELL_X1 FILLER_134_978 ();
 FILLCELL_X1 FILLER_134_1021 ();
 FILLCELL_X2 FILLER_134_1040 ();
 FILLCELL_X2 FILLER_134_1061 ();
 FILLCELL_X1 FILLER_134_1072 ();
 FILLCELL_X2 FILLER_134_1101 ();
 FILLCELL_X1 FILLER_134_1103 ();
 FILLCELL_X2 FILLER_134_1109 ();
 FILLCELL_X1 FILLER_134_1111 ();
 FILLCELL_X32 FILLER_134_1124 ();
 FILLCELL_X32 FILLER_134_1156 ();
 FILLCELL_X16 FILLER_134_1188 ();
 FILLCELL_X4 FILLER_134_1204 ();
 FILLCELL_X1 FILLER_134_1208 ();
 FILLCELL_X32 FILLER_135_1 ();
 FILLCELL_X32 FILLER_135_33 ();
 FILLCELL_X32 FILLER_135_65 ();
 FILLCELL_X32 FILLER_135_97 ();
 FILLCELL_X32 FILLER_135_129 ();
 FILLCELL_X32 FILLER_135_161 ();
 FILLCELL_X16 FILLER_135_193 ();
 FILLCELL_X8 FILLER_135_209 ();
 FILLCELL_X1 FILLER_135_243 ();
 FILLCELL_X2 FILLER_135_255 ();
 FILLCELL_X2 FILLER_135_261 ();
 FILLCELL_X4 FILLER_135_270 ();
 FILLCELL_X4 FILLER_135_283 ();
 FILLCELL_X2 FILLER_135_305 ();
 FILLCELL_X2 FILLER_135_347 ();
 FILLCELL_X1 FILLER_135_378 ();
 FILLCELL_X16 FILLER_135_391 ();
 FILLCELL_X8 FILLER_135_407 ();
 FILLCELL_X1 FILLER_135_415 ();
 FILLCELL_X2 FILLER_135_431 ();
 FILLCELL_X1 FILLER_135_433 ();
 FILLCELL_X2 FILLER_135_442 ();
 FILLCELL_X8 FILLER_135_451 ();
 FILLCELL_X1 FILLER_135_459 ();
 FILLCELL_X4 FILLER_135_467 ();
 FILLCELL_X8 FILLER_135_478 ();
 FILLCELL_X4 FILLER_135_486 ();
 FILLCELL_X4 FILLER_135_506 ();
 FILLCELL_X2 FILLER_135_513 ();
 FILLCELL_X1 FILLER_135_515 ();
 FILLCELL_X8 FILLER_135_527 ();
 FILLCELL_X2 FILLER_135_535 ();
 FILLCELL_X16 FILLER_135_546 ();
 FILLCELL_X1 FILLER_135_562 ();
 FILLCELL_X4 FILLER_135_570 ();
 FILLCELL_X4 FILLER_135_578 ();
 FILLCELL_X2 FILLER_135_600 ();
 FILLCELL_X1 FILLER_135_602 ();
 FILLCELL_X16 FILLER_135_608 ();
 FILLCELL_X8 FILLER_135_624 ();
 FILLCELL_X1 FILLER_135_632 ();
 FILLCELL_X32 FILLER_135_640 ();
 FILLCELL_X8 FILLER_135_672 ();
 FILLCELL_X2 FILLER_135_680 ();
 FILLCELL_X1 FILLER_135_682 ();
 FILLCELL_X2 FILLER_135_713 ();
 FILLCELL_X1 FILLER_135_745 ();
 FILLCELL_X1 FILLER_135_755 ();
 FILLCELL_X1 FILLER_135_780 ();
 FILLCELL_X2 FILLER_135_795 ();
 FILLCELL_X1 FILLER_135_819 ();
 FILLCELL_X1 FILLER_135_843 ();
 FILLCELL_X32 FILLER_135_851 ();
 FILLCELL_X16 FILLER_135_883 ();
 FILLCELL_X8 FILLER_135_899 ();
 FILLCELL_X4 FILLER_135_907 ();
 FILLCELL_X2 FILLER_135_911 ();
 FILLCELL_X1 FILLER_135_913 ();
 FILLCELL_X8 FILLER_135_931 ();
 FILLCELL_X2 FILLER_135_939 ();
 FILLCELL_X1 FILLER_135_950 ();
 FILLCELL_X1 FILLER_135_971 ();
 FILLCELL_X1 FILLER_135_976 ();
 FILLCELL_X1 FILLER_135_990 ();
 FILLCELL_X2 FILLER_135_1014 ();
 FILLCELL_X2 FILLER_135_1026 ();
 FILLCELL_X2 FILLER_135_1044 ();
 FILLCELL_X2 FILLER_135_1059 ();
 FILLCELL_X1 FILLER_135_1065 ();
 FILLCELL_X2 FILLER_135_1090 ();
 FILLCELL_X8 FILLER_135_1112 ();
 FILLCELL_X2 FILLER_135_1120 ();
 FILLCELL_X32 FILLER_135_1135 ();
 FILLCELL_X32 FILLER_135_1167 ();
 FILLCELL_X8 FILLER_135_1199 ();
 FILLCELL_X2 FILLER_135_1207 ();
 FILLCELL_X32 FILLER_136_1 ();
 FILLCELL_X32 FILLER_136_33 ();
 FILLCELL_X32 FILLER_136_65 ();
 FILLCELL_X32 FILLER_136_97 ();
 FILLCELL_X32 FILLER_136_129 ();
 FILLCELL_X32 FILLER_136_161 ();
 FILLCELL_X16 FILLER_136_193 ();
 FILLCELL_X4 FILLER_136_209 ();
 FILLCELL_X1 FILLER_136_213 ();
 FILLCELL_X4 FILLER_136_239 ();
 FILLCELL_X2 FILLER_136_243 ();
 FILLCELL_X2 FILLER_136_269 ();
 FILLCELL_X1 FILLER_136_271 ();
 FILLCELL_X1 FILLER_136_306 ();
 FILLCELL_X2 FILLER_136_320 ();
 FILLCELL_X1 FILLER_136_335 ();
 FILLCELL_X2 FILLER_136_347 ();
 FILLCELL_X1 FILLER_136_364 ();
 FILLCELL_X1 FILLER_136_379 ();
 FILLCELL_X8 FILLER_136_391 ();
 FILLCELL_X4 FILLER_136_399 ();
 FILLCELL_X2 FILLER_136_403 ();
 FILLCELL_X1 FILLER_136_405 ();
 FILLCELL_X16 FILLER_136_423 ();
 FILLCELL_X8 FILLER_136_439 ();
 FILLCELL_X4 FILLER_136_447 ();
 FILLCELL_X2 FILLER_136_451 ();
 FILLCELL_X1 FILLER_136_456 ();
 FILLCELL_X1 FILLER_136_461 ();
 FILLCELL_X1 FILLER_136_470 ();
 FILLCELL_X2 FILLER_136_479 ();
 FILLCELL_X1 FILLER_136_481 ();
 FILLCELL_X8 FILLER_136_494 ();
 FILLCELL_X4 FILLER_136_502 ();
 FILLCELL_X1 FILLER_136_506 ();
 FILLCELL_X4 FILLER_136_515 ();
 FILLCELL_X2 FILLER_136_533 ();
 FILLCELL_X4 FILLER_136_539 ();
 FILLCELL_X4 FILLER_136_548 ();
 FILLCELL_X2 FILLER_136_571 ();
 FILLCELL_X2 FILLER_136_584 ();
 FILLCELL_X1 FILLER_136_586 ();
 FILLCELL_X8 FILLER_136_592 ();
 FILLCELL_X4 FILLER_136_609 ();
 FILLCELL_X1 FILLER_136_613 ();
 FILLCELL_X16 FILLER_136_632 ();
 FILLCELL_X8 FILLER_136_648 ();
 FILLCELL_X2 FILLER_136_656 ();
 FILLCELL_X1 FILLER_136_658 ();
 FILLCELL_X4 FILLER_136_677 ();
 FILLCELL_X4 FILLER_136_694 ();
 FILLCELL_X2 FILLER_136_698 ();
 FILLCELL_X1 FILLER_136_700 ();
 FILLCELL_X2 FILLER_136_710 ();
 FILLCELL_X1 FILLER_136_712 ();
 FILLCELL_X4 FILLER_136_716 ();
 FILLCELL_X2 FILLER_136_720 ();
 FILLCELL_X1 FILLER_136_722 ();
 FILLCELL_X1 FILLER_136_726 ();
 FILLCELL_X1 FILLER_136_739 ();
 FILLCELL_X4 FILLER_136_777 ();
 FILLCELL_X1 FILLER_136_781 ();
 FILLCELL_X4 FILLER_136_789 ();
 FILLCELL_X2 FILLER_136_797 ();
 FILLCELL_X1 FILLER_136_799 ();
 FILLCELL_X4 FILLER_136_813 ();
 FILLCELL_X1 FILLER_136_822 ();
 FILLCELL_X8 FILLER_136_838 ();
 FILLCELL_X4 FILLER_136_846 ();
 FILLCELL_X2 FILLER_136_850 ();
 FILLCELL_X1 FILLER_136_852 ();
 FILLCELL_X32 FILLER_136_860 ();
 FILLCELL_X2 FILLER_136_892 ();
 FILLCELL_X32 FILLER_136_901 ();
 FILLCELL_X2 FILLER_136_933 ();
 FILLCELL_X2 FILLER_136_951 ();
 FILLCELL_X1 FILLER_136_968 ();
 FILLCELL_X1 FILLER_136_991 ();
 FILLCELL_X8 FILLER_136_1078 ();
 FILLCELL_X2 FILLER_136_1086 ();
 FILLCELL_X2 FILLER_136_1092 ();
 FILLCELL_X1 FILLER_136_1094 ();
 FILLCELL_X2 FILLER_136_1098 ();
 FILLCELL_X4 FILLER_136_1106 ();
 FILLCELL_X2 FILLER_136_1113 ();
 FILLCELL_X1 FILLER_136_1115 ();
 FILLCELL_X8 FILLER_136_1125 ();
 FILLCELL_X2 FILLER_136_1133 ();
 FILLCELL_X32 FILLER_136_1138 ();
 FILLCELL_X32 FILLER_136_1170 ();
 FILLCELL_X4 FILLER_136_1202 ();
 FILLCELL_X2 FILLER_136_1206 ();
 FILLCELL_X1 FILLER_136_1208 ();
 FILLCELL_X32 FILLER_137_1 ();
 FILLCELL_X32 FILLER_137_33 ();
 FILLCELL_X32 FILLER_137_65 ();
 FILLCELL_X32 FILLER_137_97 ();
 FILLCELL_X32 FILLER_137_129 ();
 FILLCELL_X32 FILLER_137_161 ();
 FILLCELL_X32 FILLER_137_193 ();
 FILLCELL_X2 FILLER_137_225 ();
 FILLCELL_X1 FILLER_137_227 ();
 FILLCELL_X4 FILLER_137_235 ();
 FILLCELL_X2 FILLER_137_239 ();
 FILLCELL_X8 FILLER_137_244 ();
 FILLCELL_X4 FILLER_137_252 ();
 FILLCELL_X4 FILLER_137_281 ();
 FILLCELL_X2 FILLER_137_285 ();
 FILLCELL_X1 FILLER_137_287 ();
 FILLCELL_X1 FILLER_137_314 ();
 FILLCELL_X1 FILLER_137_350 ();
 FILLCELL_X2 FILLER_137_356 ();
 FILLCELL_X2 FILLER_137_362 ();
 FILLCELL_X2 FILLER_137_375 ();
 FILLCELL_X1 FILLER_137_377 ();
 FILLCELL_X16 FILLER_137_394 ();
 FILLCELL_X8 FILLER_137_410 ();
 FILLCELL_X4 FILLER_137_418 ();
 FILLCELL_X4 FILLER_137_439 ();
 FILLCELL_X2 FILLER_137_443 ();
 FILLCELL_X1 FILLER_137_452 ();
 FILLCELL_X1 FILLER_137_457 ();
 FILLCELL_X2 FILLER_137_466 ();
 FILLCELL_X1 FILLER_137_475 ();
 FILLCELL_X4 FILLER_137_495 ();
 FILLCELL_X2 FILLER_137_499 ();
 FILLCELL_X1 FILLER_137_501 ();
 FILLCELL_X8 FILLER_137_525 ();
 FILLCELL_X1 FILLER_137_533 ();
 FILLCELL_X4 FILLER_137_540 ();
 FILLCELL_X2 FILLER_137_544 ();
 FILLCELL_X1 FILLER_137_550 ();
 FILLCELL_X1 FILLER_137_555 ();
 FILLCELL_X4 FILLER_137_578 ();
 FILLCELL_X2 FILLER_137_582 ();
 FILLCELL_X32 FILLER_137_598 ();
 FILLCELL_X32 FILLER_137_630 ();
 FILLCELL_X8 FILLER_137_662 ();
 FILLCELL_X1 FILLER_137_670 ();
 FILLCELL_X4 FILLER_137_684 ();
 FILLCELL_X2 FILLER_137_688 ();
 FILLCELL_X2 FILLER_137_700 ();
 FILLCELL_X2 FILLER_137_706 ();
 FILLCELL_X1 FILLER_137_708 ();
 FILLCELL_X1 FILLER_137_712 ();
 FILLCELL_X8 FILLER_137_779 ();
 FILLCELL_X2 FILLER_137_787 ();
 FILLCELL_X2 FILLER_137_809 ();
 FILLCELL_X1 FILLER_137_811 ();
 FILLCELL_X2 FILLER_137_845 ();
 FILLCELL_X1 FILLER_137_847 ();
 FILLCELL_X32 FILLER_137_874 ();
 FILLCELL_X4 FILLER_137_906 ();
 FILLCELL_X8 FILLER_137_929 ();
 FILLCELL_X1 FILLER_137_937 ();
 FILLCELL_X2 FILLER_137_998 ();
 FILLCELL_X2 FILLER_137_1038 ();
 FILLCELL_X4 FILLER_137_1076 ();
 FILLCELL_X2 FILLER_137_1080 ();
 FILLCELL_X2 FILLER_137_1087 ();
 FILLCELL_X1 FILLER_137_1092 ();
 FILLCELL_X2 FILLER_137_1104 ();
 FILLCELL_X1 FILLER_137_1106 ();
 FILLCELL_X2 FILLER_137_1121 ();
 FILLCELL_X32 FILLER_137_1127 ();
 FILLCELL_X32 FILLER_137_1159 ();
 FILLCELL_X16 FILLER_137_1191 ();
 FILLCELL_X2 FILLER_137_1207 ();
 FILLCELL_X32 FILLER_138_1 ();
 FILLCELL_X32 FILLER_138_33 ();
 FILLCELL_X32 FILLER_138_65 ();
 FILLCELL_X32 FILLER_138_97 ();
 FILLCELL_X32 FILLER_138_129 ();
 FILLCELL_X32 FILLER_138_161 ();
 FILLCELL_X16 FILLER_138_193 ();
 FILLCELL_X2 FILLER_138_209 ();
 FILLCELL_X4 FILLER_138_224 ();
 FILLCELL_X1 FILLER_138_228 ();
 FILLCELL_X2 FILLER_138_232 ();
 FILLCELL_X1 FILLER_138_234 ();
 FILLCELL_X4 FILLER_138_263 ();
 FILLCELL_X1 FILLER_138_267 ();
 FILLCELL_X1 FILLER_138_272 ();
 FILLCELL_X1 FILLER_138_283 ();
 FILLCELL_X2 FILLER_138_292 ();
 FILLCELL_X1 FILLER_138_306 ();
 FILLCELL_X4 FILLER_138_314 ();
 FILLCELL_X1 FILLER_138_329 ();
 FILLCELL_X1 FILLER_138_334 ();
 FILLCELL_X4 FILLER_138_344 ();
 FILLCELL_X1 FILLER_138_348 ();
 FILLCELL_X2 FILLER_138_362 ();
 FILLCELL_X1 FILLER_138_371 ();
 FILLCELL_X1 FILLER_138_376 ();
 FILLCELL_X8 FILLER_138_388 ();
 FILLCELL_X4 FILLER_138_396 ();
 FILLCELL_X16 FILLER_138_407 ();
 FILLCELL_X8 FILLER_138_423 ();
 FILLCELL_X2 FILLER_138_431 ();
 FILLCELL_X1 FILLER_138_433 ();
 FILLCELL_X2 FILLER_138_471 ();
 FILLCELL_X1 FILLER_138_473 ();
 FILLCELL_X4 FILLER_138_490 ();
 FILLCELL_X1 FILLER_138_494 ();
 FILLCELL_X4 FILLER_138_499 ();
 FILLCELL_X2 FILLER_138_541 ();
 FILLCELL_X2 FILLER_138_562 ();
 FILLCELL_X1 FILLER_138_564 ();
 FILLCELL_X4 FILLER_138_572 ();
 FILLCELL_X1 FILLER_138_576 ();
 FILLCELL_X8 FILLER_138_621 ();
 FILLCELL_X2 FILLER_138_629 ();
 FILLCELL_X32 FILLER_138_632 ();
 FILLCELL_X8 FILLER_138_664 ();
 FILLCELL_X2 FILLER_138_672 ();
 FILLCELL_X2 FILLER_138_700 ();
 FILLCELL_X2 FILLER_138_713 ();
 FILLCELL_X2 FILLER_138_734 ();
 FILLCELL_X1 FILLER_138_743 ();
 FILLCELL_X2 FILLER_138_758 ();
 FILLCELL_X1 FILLER_138_760 ();
 FILLCELL_X8 FILLER_138_776 ();
 FILLCELL_X2 FILLER_138_788 ();
 FILLCELL_X8 FILLER_138_811 ();
 FILLCELL_X2 FILLER_138_819 ();
 FILLCELL_X1 FILLER_138_821 ();
 FILLCELL_X1 FILLER_138_826 ();
 FILLCELL_X1 FILLER_138_840 ();
 FILLCELL_X2 FILLER_138_852 ();
 FILLCELL_X8 FILLER_138_870 ();
 FILLCELL_X32 FILLER_138_895 ();
 FILLCELL_X8 FILLER_138_927 ();
 FILLCELL_X1 FILLER_138_935 ();
 FILLCELL_X1 FILLER_138_973 ();
 FILLCELL_X1 FILLER_138_1014 ();
 FILLCELL_X2 FILLER_138_1030 ();
 FILLCELL_X2 FILLER_138_1048 ();
 FILLCELL_X1 FILLER_138_1059 ();
 FILLCELL_X2 FILLER_138_1071 ();
 FILLCELL_X1 FILLER_138_1115 ();
 FILLCELL_X32 FILLER_138_1141 ();
 FILLCELL_X32 FILLER_138_1173 ();
 FILLCELL_X4 FILLER_138_1205 ();
 FILLCELL_X32 FILLER_139_1 ();
 FILLCELL_X32 FILLER_139_33 ();
 FILLCELL_X32 FILLER_139_65 ();
 FILLCELL_X32 FILLER_139_97 ();
 FILLCELL_X32 FILLER_139_129 ();
 FILLCELL_X32 FILLER_139_161 ();
 FILLCELL_X16 FILLER_139_193 ();
 FILLCELL_X8 FILLER_139_209 ();
 FILLCELL_X4 FILLER_139_217 ();
 FILLCELL_X2 FILLER_139_245 ();
 FILLCELL_X1 FILLER_139_247 ();
 FILLCELL_X2 FILLER_139_255 ();
 FILLCELL_X1 FILLER_139_290 ();
 FILLCELL_X16 FILLER_139_314 ();
 FILLCELL_X4 FILLER_139_330 ();
 FILLCELL_X2 FILLER_139_334 ();
 FILLCELL_X1 FILLER_139_336 ();
 FILLCELL_X1 FILLER_139_340 ();
 FILLCELL_X1 FILLER_139_375 ();
 FILLCELL_X2 FILLER_139_397 ();
 FILLCELL_X32 FILLER_139_410 ();
 FILLCELL_X8 FILLER_139_442 ();
 FILLCELL_X2 FILLER_139_450 ();
 FILLCELL_X1 FILLER_139_452 ();
 FILLCELL_X8 FILLER_139_462 ();
 FILLCELL_X4 FILLER_139_480 ();
 FILLCELL_X8 FILLER_139_492 ();
 FILLCELL_X1 FILLER_139_500 ();
 FILLCELL_X16 FILLER_139_509 ();
 FILLCELL_X2 FILLER_139_529 ();
 FILLCELL_X1 FILLER_139_531 ();
 FILLCELL_X16 FILLER_139_543 ();
 FILLCELL_X4 FILLER_139_559 ();
 FILLCELL_X1 FILLER_139_563 ();
 FILLCELL_X16 FILLER_139_600 ();
 FILLCELL_X1 FILLER_139_616 ();
 FILLCELL_X16 FILLER_139_639 ();
 FILLCELL_X4 FILLER_139_655 ();
 FILLCELL_X8 FILLER_139_672 ();
 FILLCELL_X2 FILLER_139_680 ();
 FILLCELL_X1 FILLER_139_682 ();
 FILLCELL_X2 FILLER_139_735 ();
 FILLCELL_X1 FILLER_139_737 ();
 FILLCELL_X2 FILLER_139_741 ();
 FILLCELL_X1 FILLER_139_743 ();
 FILLCELL_X8 FILLER_139_754 ();
 FILLCELL_X2 FILLER_139_769 ();
 FILLCELL_X1 FILLER_139_771 ();
 FILLCELL_X2 FILLER_139_775 ();
 FILLCELL_X1 FILLER_139_777 ();
 FILLCELL_X1 FILLER_139_798 ();
 FILLCELL_X2 FILLER_139_832 ();
 FILLCELL_X4 FILLER_139_844 ();
 FILLCELL_X4 FILLER_139_853 ();
 FILLCELL_X2 FILLER_139_878 ();
 FILLCELL_X4 FILLER_139_887 ();
 FILLCELL_X2 FILLER_139_891 ();
 FILLCELL_X16 FILLER_139_910 ();
 FILLCELL_X8 FILLER_139_926 ();
 FILLCELL_X1 FILLER_139_934 ();
 FILLCELL_X2 FILLER_139_948 ();
 FILLCELL_X2 FILLER_139_953 ();
 FILLCELL_X1 FILLER_139_955 ();
 FILLCELL_X1 FILLER_139_992 ();
 FILLCELL_X1 FILLER_139_1029 ();
 FILLCELL_X2 FILLER_139_1039 ();
 FILLCELL_X1 FILLER_139_1060 ();
 FILLCELL_X2 FILLER_139_1073 ();
 FILLCELL_X1 FILLER_139_1090 ();
 FILLCELL_X32 FILLER_139_1132 ();
 FILLCELL_X32 FILLER_139_1164 ();
 FILLCELL_X8 FILLER_139_1196 ();
 FILLCELL_X4 FILLER_139_1204 ();
 FILLCELL_X1 FILLER_139_1208 ();
 FILLCELL_X32 FILLER_140_1 ();
 FILLCELL_X32 FILLER_140_33 ();
 FILLCELL_X32 FILLER_140_65 ();
 FILLCELL_X32 FILLER_140_97 ();
 FILLCELL_X32 FILLER_140_129 ();
 FILLCELL_X32 FILLER_140_161 ();
 FILLCELL_X32 FILLER_140_193 ();
 FILLCELL_X4 FILLER_140_225 ();
 FILLCELL_X1 FILLER_140_229 ();
 FILLCELL_X4 FILLER_140_247 ();
 FILLCELL_X1 FILLER_140_251 ();
 FILLCELL_X1 FILLER_140_265 ();
 FILLCELL_X1 FILLER_140_285 ();
 FILLCELL_X2 FILLER_140_296 ();
 FILLCELL_X4 FILLER_140_314 ();
 FILLCELL_X1 FILLER_140_318 ();
 FILLCELL_X4 FILLER_140_328 ();
 FILLCELL_X2 FILLER_140_332 ();
 FILLCELL_X4 FILLER_140_353 ();
 FILLCELL_X2 FILLER_140_359 ();
 FILLCELL_X4 FILLER_140_364 ();
 FILLCELL_X2 FILLER_140_368 ();
 FILLCELL_X4 FILLER_140_375 ();
 FILLCELL_X32 FILLER_140_396 ();
 FILLCELL_X16 FILLER_140_428 ();
 FILLCELL_X8 FILLER_140_444 ();
 FILLCELL_X4 FILLER_140_452 ();
 FILLCELL_X2 FILLER_140_456 ();
 FILLCELL_X1 FILLER_140_458 ();
 FILLCELL_X1 FILLER_140_479 ();
 FILLCELL_X2 FILLER_140_484 ();
 FILLCELL_X4 FILLER_140_492 ();
 FILLCELL_X2 FILLER_140_496 ();
 FILLCELL_X1 FILLER_140_500 ();
 FILLCELL_X4 FILLER_140_513 ();
 FILLCELL_X1 FILLER_140_517 ();
 FILLCELL_X16 FILLER_140_525 ();
 FILLCELL_X1 FILLER_140_541 ();
 FILLCELL_X4 FILLER_140_554 ();
 FILLCELL_X1 FILLER_140_565 ();
 FILLCELL_X2 FILLER_140_575 ();
 FILLCELL_X2 FILLER_140_586 ();
 FILLCELL_X1 FILLER_140_592 ();
 FILLCELL_X1 FILLER_140_609 ();
 FILLCELL_X4 FILLER_140_613 ();
 FILLCELL_X2 FILLER_140_629 ();
 FILLCELL_X32 FILLER_140_632 ();
 FILLCELL_X8 FILLER_140_664 ();
 FILLCELL_X4 FILLER_140_672 ();
 FILLCELL_X2 FILLER_140_685 ();
 FILLCELL_X2 FILLER_140_696 ();
 FILLCELL_X4 FILLER_140_703 ();
 FILLCELL_X2 FILLER_140_707 ();
 FILLCELL_X1 FILLER_140_709 ();
 FILLCELL_X1 FILLER_140_729 ();
 FILLCELL_X2 FILLER_140_749 ();
 FILLCELL_X2 FILLER_140_756 ();
 FILLCELL_X1 FILLER_140_758 ();
 FILLCELL_X1 FILLER_140_762 ();
 FILLCELL_X2 FILLER_140_776 ();
 FILLCELL_X2 FILLER_140_784 ();
 FILLCELL_X4 FILLER_140_797 ();
 FILLCELL_X4 FILLER_140_817 ();
 FILLCELL_X1 FILLER_140_821 ();
 FILLCELL_X1 FILLER_140_840 ();
 FILLCELL_X1 FILLER_140_850 ();
 FILLCELL_X1 FILLER_140_858 ();
 FILLCELL_X32 FILLER_140_878 ();
 FILLCELL_X32 FILLER_140_910 ();
 FILLCELL_X2 FILLER_140_942 ();
 FILLCELL_X1 FILLER_140_957 ();
 FILLCELL_X1 FILLER_140_983 ();
 FILLCELL_X1 FILLER_140_993 ();
 FILLCELL_X1 FILLER_140_1011 ();
 FILLCELL_X2 FILLER_140_1021 ();
 FILLCELL_X1 FILLER_140_1023 ();
 FILLCELL_X2 FILLER_140_1031 ();
 FILLCELL_X2 FILLER_140_1055 ();
 FILLCELL_X4 FILLER_140_1062 ();
 FILLCELL_X2 FILLER_140_1066 ();
 FILLCELL_X1 FILLER_140_1068 ();
 FILLCELL_X1 FILLER_140_1123 ();
 FILLCELL_X4 FILLER_140_1133 ();
 FILLCELL_X32 FILLER_140_1147 ();
 FILLCELL_X16 FILLER_140_1179 ();
 FILLCELL_X8 FILLER_140_1195 ();
 FILLCELL_X4 FILLER_140_1203 ();
 FILLCELL_X2 FILLER_140_1207 ();
 FILLCELL_X32 FILLER_141_1 ();
 FILLCELL_X32 FILLER_141_33 ();
 FILLCELL_X32 FILLER_141_65 ();
 FILLCELL_X32 FILLER_141_97 ();
 FILLCELL_X32 FILLER_141_129 ();
 FILLCELL_X32 FILLER_141_161 ();
 FILLCELL_X16 FILLER_141_193 ();
 FILLCELL_X8 FILLER_141_209 ();
 FILLCELL_X4 FILLER_141_217 ();
 FILLCELL_X2 FILLER_141_221 ();
 FILLCELL_X1 FILLER_141_223 ();
 FILLCELL_X1 FILLER_141_279 ();
 FILLCELL_X2 FILLER_141_302 ();
 FILLCELL_X1 FILLER_141_304 ();
 FILLCELL_X2 FILLER_141_309 ();
 FILLCELL_X1 FILLER_141_311 ();
 FILLCELL_X8 FILLER_141_319 ();
 FILLCELL_X2 FILLER_141_327 ();
 FILLCELL_X4 FILLER_141_340 ();
 FILLCELL_X1 FILLER_141_344 ();
 FILLCELL_X1 FILLER_141_360 ();
 FILLCELL_X1 FILLER_141_383 ();
 FILLCELL_X32 FILLER_141_401 ();
 FILLCELL_X8 FILLER_141_433 ();
 FILLCELL_X4 FILLER_141_441 ();
 FILLCELL_X2 FILLER_141_445 ();
 FILLCELL_X1 FILLER_141_447 ();
 FILLCELL_X2 FILLER_141_484 ();
 FILLCELL_X1 FILLER_141_486 ();
 FILLCELL_X1 FILLER_141_495 ();
 FILLCELL_X4 FILLER_141_516 ();
 FILLCELL_X2 FILLER_141_528 ();
 FILLCELL_X1 FILLER_141_530 ();
 FILLCELL_X2 FILLER_141_541 ();
 FILLCELL_X1 FILLER_141_543 ();
 FILLCELL_X4 FILLER_141_555 ();
 FILLCELL_X2 FILLER_141_564 ();
 FILLCELL_X1 FILLER_141_566 ();
 FILLCELL_X2 FILLER_141_574 ();
 FILLCELL_X1 FILLER_141_576 ();
 FILLCELL_X1 FILLER_141_594 ();
 FILLCELL_X32 FILLER_141_620 ();
 FILLCELL_X16 FILLER_141_652 ();
 FILLCELL_X8 FILLER_141_668 ();
 FILLCELL_X4 FILLER_141_676 ();
 FILLCELL_X1 FILLER_141_680 ();
 FILLCELL_X2 FILLER_141_701 ();
 FILLCELL_X1 FILLER_141_703 ();
 FILLCELL_X1 FILLER_141_711 ();
 FILLCELL_X2 FILLER_141_742 ();
 FILLCELL_X1 FILLER_141_744 ();
 FILLCELL_X1 FILLER_141_756 ();
 FILLCELL_X1 FILLER_141_775 ();
 FILLCELL_X8 FILLER_141_787 ();
 FILLCELL_X4 FILLER_141_795 ();
 FILLCELL_X1 FILLER_141_799 ();
 FILLCELL_X2 FILLER_141_805 ();
 FILLCELL_X1 FILLER_141_811 ();
 FILLCELL_X1 FILLER_141_816 ();
 FILLCELL_X2 FILLER_141_822 ();
 FILLCELL_X1 FILLER_141_824 ();
 FILLCELL_X2 FILLER_141_845 ();
 FILLCELL_X1 FILLER_141_847 ();
 FILLCELL_X2 FILLER_141_853 ();
 FILLCELL_X1 FILLER_141_866 ();
 FILLCELL_X4 FILLER_141_873 ();
 FILLCELL_X8 FILLER_141_883 ();
 FILLCELL_X4 FILLER_141_891 ();
 FILLCELL_X2 FILLER_141_895 ();
 FILLCELL_X16 FILLER_141_914 ();
 FILLCELL_X8 FILLER_141_930 ();
 FILLCELL_X2 FILLER_141_938 ();
 FILLCELL_X1 FILLER_141_940 ();
 FILLCELL_X4 FILLER_141_959 ();
 FILLCELL_X2 FILLER_141_966 ();
 FILLCELL_X1 FILLER_141_990 ();
 FILLCELL_X2 FILLER_141_996 ();
 FILLCELL_X2 FILLER_141_1005 ();
 FILLCELL_X1 FILLER_141_1007 ();
 FILLCELL_X1 FILLER_141_1017 ();
 FILLCELL_X1 FILLER_141_1042 ();
 FILLCELL_X1 FILLER_141_1051 ();
 FILLCELL_X2 FILLER_141_1070 ();
 FILLCELL_X1 FILLER_141_1072 ();
 FILLCELL_X1 FILLER_141_1078 ();
 FILLCELL_X2 FILLER_141_1086 ();
 FILLCELL_X32 FILLER_141_1132 ();
 FILLCELL_X32 FILLER_141_1164 ();
 FILLCELL_X8 FILLER_141_1196 ();
 FILLCELL_X4 FILLER_141_1204 ();
 FILLCELL_X1 FILLER_141_1208 ();
 FILLCELL_X32 FILLER_142_1 ();
 FILLCELL_X32 FILLER_142_33 ();
 FILLCELL_X32 FILLER_142_65 ();
 FILLCELL_X32 FILLER_142_97 ();
 FILLCELL_X32 FILLER_142_129 ();
 FILLCELL_X32 FILLER_142_161 ();
 FILLCELL_X16 FILLER_142_193 ();
 FILLCELL_X1 FILLER_142_209 ();
 FILLCELL_X16 FILLER_142_281 ();
 FILLCELL_X1 FILLER_142_297 ();
 FILLCELL_X2 FILLER_142_300 ();
 FILLCELL_X2 FILLER_142_323 ();
 FILLCELL_X1 FILLER_142_325 ();
 FILLCELL_X4 FILLER_142_330 ();
 FILLCELL_X2 FILLER_142_334 ();
 FILLCELL_X2 FILLER_142_347 ();
 FILLCELL_X1 FILLER_142_349 ();
 FILLCELL_X1 FILLER_142_364 ();
 FILLCELL_X4 FILLER_142_376 ();
 FILLCELL_X2 FILLER_142_380 ();
 FILLCELL_X1 FILLER_142_382 ();
 FILLCELL_X1 FILLER_142_399 ();
 FILLCELL_X32 FILLER_142_405 ();
 FILLCELL_X8 FILLER_142_437 ();
 FILLCELL_X4 FILLER_142_445 ();
 FILLCELL_X2 FILLER_142_449 ();
 FILLCELL_X1 FILLER_142_451 ();
 FILLCELL_X2 FILLER_142_469 ();
 FILLCELL_X4 FILLER_142_490 ();
 FILLCELL_X1 FILLER_142_494 ();
 FILLCELL_X4 FILLER_142_501 ();
 FILLCELL_X2 FILLER_142_505 ();
 FILLCELL_X1 FILLER_142_507 ();
 FILLCELL_X8 FILLER_142_512 ();
 FILLCELL_X1 FILLER_142_520 ();
 FILLCELL_X8 FILLER_142_529 ();
 FILLCELL_X4 FILLER_142_537 ();
 FILLCELL_X1 FILLER_142_541 ();
 FILLCELL_X1 FILLER_142_546 ();
 FILLCELL_X2 FILLER_142_558 ();
 FILLCELL_X1 FILLER_142_564 ();
 FILLCELL_X2 FILLER_142_576 ();
 FILLCELL_X8 FILLER_142_619 ();
 FILLCELL_X4 FILLER_142_627 ();
 FILLCELL_X32 FILLER_142_632 ();
 FILLCELL_X8 FILLER_142_664 ();
 FILLCELL_X4 FILLER_142_672 ();
 FILLCELL_X1 FILLER_142_676 ();
 FILLCELL_X1 FILLER_142_690 ();
 FILLCELL_X4 FILLER_142_700 ();
 FILLCELL_X1 FILLER_142_722 ();
 FILLCELL_X4 FILLER_142_756 ();
 FILLCELL_X8 FILLER_142_773 ();
 FILLCELL_X1 FILLER_142_785 ();
 FILLCELL_X1 FILLER_142_790 ();
 FILLCELL_X4 FILLER_142_795 ();
 FILLCELL_X1 FILLER_142_799 ();
 FILLCELL_X2 FILLER_142_804 ();
 FILLCELL_X1 FILLER_142_806 ();
 FILLCELL_X8 FILLER_142_813 ();
 FILLCELL_X1 FILLER_142_837 ();
 FILLCELL_X1 FILLER_142_842 ();
 FILLCELL_X1 FILLER_142_847 ();
 FILLCELL_X1 FILLER_142_851 ();
 FILLCELL_X2 FILLER_142_855 ();
 FILLCELL_X1 FILLER_142_857 ();
 FILLCELL_X1 FILLER_142_868 ();
 FILLCELL_X4 FILLER_142_873 ();
 FILLCELL_X2 FILLER_142_877 ();
 FILLCELL_X16 FILLER_142_886 ();
 FILLCELL_X8 FILLER_142_902 ();
 FILLCELL_X4 FILLER_142_910 ();
 FILLCELL_X2 FILLER_142_914 ();
 FILLCELL_X1 FILLER_142_916 ();
 FILLCELL_X8 FILLER_142_925 ();
 FILLCELL_X2 FILLER_142_933 ();
 FILLCELL_X1 FILLER_142_1014 ();
 FILLCELL_X2 FILLER_142_1040 ();
 FILLCELL_X8 FILLER_142_1056 ();
 FILLCELL_X2 FILLER_142_1064 ();
 FILLCELL_X2 FILLER_142_1070 ();
 FILLCELL_X1 FILLER_142_1076 ();
 FILLCELL_X4 FILLER_142_1083 ();
 FILLCELL_X2 FILLER_142_1087 ();
 FILLCELL_X4 FILLER_142_1121 ();
 FILLCELL_X2 FILLER_142_1127 ();
 FILLCELL_X1 FILLER_142_1129 ();
 FILLCELL_X32 FILLER_142_1133 ();
 FILLCELL_X32 FILLER_142_1165 ();
 FILLCELL_X8 FILLER_142_1197 ();
 FILLCELL_X4 FILLER_142_1205 ();
 FILLCELL_X32 FILLER_143_1 ();
 FILLCELL_X32 FILLER_143_33 ();
 FILLCELL_X32 FILLER_143_65 ();
 FILLCELL_X32 FILLER_143_97 ();
 FILLCELL_X32 FILLER_143_129 ();
 FILLCELL_X32 FILLER_143_161 ();
 FILLCELL_X16 FILLER_143_193 ();
 FILLCELL_X2 FILLER_143_209 ();
 FILLCELL_X1 FILLER_143_211 ();
 FILLCELL_X1 FILLER_143_253 ();
 FILLCELL_X1 FILLER_143_258 ();
 FILLCELL_X2 FILLER_143_283 ();
 FILLCELL_X1 FILLER_143_289 ();
 FILLCELL_X2 FILLER_143_294 ();
 FILLCELL_X4 FILLER_143_303 ();
 FILLCELL_X1 FILLER_143_332 ();
 FILLCELL_X1 FILLER_143_339 ();
 FILLCELL_X1 FILLER_143_351 ();
 FILLCELL_X8 FILLER_143_363 ();
 FILLCELL_X2 FILLER_143_375 ();
 FILLCELL_X1 FILLER_143_377 ();
 FILLCELL_X4 FILLER_143_382 ();
 FILLCELL_X1 FILLER_143_386 ();
 FILLCELL_X32 FILLER_143_404 ();
 FILLCELL_X8 FILLER_143_436 ();
 FILLCELL_X4 FILLER_143_444 ();
 FILLCELL_X2 FILLER_143_466 ();
 FILLCELL_X1 FILLER_143_468 ();
 FILLCELL_X2 FILLER_143_477 ();
 FILLCELL_X1 FILLER_143_479 ();
 FILLCELL_X8 FILLER_143_494 ();
 FILLCELL_X4 FILLER_143_502 ();
 FILLCELL_X2 FILLER_143_516 ();
 FILLCELL_X2 FILLER_143_525 ();
 FILLCELL_X2 FILLER_143_531 ();
 FILLCELL_X8 FILLER_143_541 ();
 FILLCELL_X1 FILLER_143_549 ();
 FILLCELL_X1 FILLER_143_561 ();
 FILLCELL_X1 FILLER_143_566 ();
 FILLCELL_X1 FILLER_143_574 ();
 FILLCELL_X32 FILLER_143_614 ();
 FILLCELL_X32 FILLER_143_646 ();
 FILLCELL_X1 FILLER_143_678 ();
 FILLCELL_X2 FILLER_143_686 ();
 FILLCELL_X1 FILLER_143_688 ();
 FILLCELL_X2 FILLER_143_702 ();
 FILLCELL_X1 FILLER_143_704 ();
 FILLCELL_X1 FILLER_143_727 ();
 FILLCELL_X8 FILLER_143_738 ();
 FILLCELL_X4 FILLER_143_746 ();
 FILLCELL_X2 FILLER_143_750 ();
 FILLCELL_X1 FILLER_143_752 ();
 FILLCELL_X8 FILLER_143_760 ();
 FILLCELL_X1 FILLER_143_771 ();
 FILLCELL_X2 FILLER_143_775 ();
 FILLCELL_X1 FILLER_143_777 ();
 FILLCELL_X4 FILLER_143_791 ();
 FILLCELL_X2 FILLER_143_795 ();
 FILLCELL_X1 FILLER_143_797 ();
 FILLCELL_X4 FILLER_143_811 ();
 FILLCELL_X1 FILLER_143_815 ();
 FILLCELL_X4 FILLER_143_819 ();
 FILLCELL_X2 FILLER_143_823 ();
 FILLCELL_X1 FILLER_143_835 ();
 FILLCELL_X4 FILLER_143_865 ();
 FILLCELL_X2 FILLER_143_869 ();
 FILLCELL_X1 FILLER_143_879 ();
 FILLCELL_X32 FILLER_143_882 ();
 FILLCELL_X16 FILLER_143_914 ();
 FILLCELL_X2 FILLER_143_930 ();
 FILLCELL_X1 FILLER_143_932 ();
 FILLCELL_X1 FILLER_143_971 ();
 FILLCELL_X2 FILLER_143_983 ();
 FILLCELL_X1 FILLER_143_1011 ();
 FILLCELL_X4 FILLER_143_1044 ();
 FILLCELL_X2 FILLER_143_1048 ();
 FILLCELL_X1 FILLER_143_1050 ();
 FILLCELL_X4 FILLER_143_1072 ();
 FILLCELL_X4 FILLER_143_1098 ();
 FILLCELL_X1 FILLER_143_1102 ();
 FILLCELL_X1 FILLER_143_1107 ();
 FILLCELL_X2 FILLER_143_1131 ();
 FILLCELL_X32 FILLER_143_1144 ();
 FILLCELL_X32 FILLER_143_1176 ();
 FILLCELL_X1 FILLER_143_1208 ();
 FILLCELL_X32 FILLER_144_1 ();
 FILLCELL_X32 FILLER_144_33 ();
 FILLCELL_X32 FILLER_144_65 ();
 FILLCELL_X32 FILLER_144_97 ();
 FILLCELL_X32 FILLER_144_129 ();
 FILLCELL_X32 FILLER_144_161 ();
 FILLCELL_X4 FILLER_144_193 ();
 FILLCELL_X1 FILLER_144_197 ();
 FILLCELL_X1 FILLER_144_230 ();
 FILLCELL_X2 FILLER_144_235 ();
 FILLCELL_X2 FILLER_144_247 ();
 FILLCELL_X1 FILLER_144_259 ();
 FILLCELL_X16 FILLER_144_288 ();
 FILLCELL_X8 FILLER_144_304 ();
 FILLCELL_X4 FILLER_144_312 ();
 FILLCELL_X2 FILLER_144_316 ();
 FILLCELL_X1 FILLER_144_318 ();
 FILLCELL_X8 FILLER_144_330 ();
 FILLCELL_X2 FILLER_144_338 ();
 FILLCELL_X1 FILLER_144_340 ();
 FILLCELL_X4 FILLER_144_345 ();
 FILLCELL_X4 FILLER_144_355 ();
 FILLCELL_X1 FILLER_144_359 ();
 FILLCELL_X1 FILLER_144_363 ();
 FILLCELL_X1 FILLER_144_378 ();
 FILLCELL_X4 FILLER_144_383 ();
 FILLCELL_X1 FILLER_144_387 ();
 FILLCELL_X1 FILLER_144_391 ();
 FILLCELL_X32 FILLER_144_400 ();
 FILLCELL_X8 FILLER_144_432 ();
 FILLCELL_X4 FILLER_144_440 ();
 FILLCELL_X2 FILLER_144_444 ();
 FILLCELL_X1 FILLER_144_446 ();
 FILLCELL_X2 FILLER_144_450 ();
 FILLCELL_X1 FILLER_144_462 ();
 FILLCELL_X2 FILLER_144_479 ();
 FILLCELL_X4 FILLER_144_485 ();
 FILLCELL_X2 FILLER_144_489 ();
 FILLCELL_X1 FILLER_144_491 ();
 FILLCELL_X8 FILLER_144_510 ();
 FILLCELL_X16 FILLER_144_525 ();
 FILLCELL_X8 FILLER_144_541 ();
 FILLCELL_X4 FILLER_144_549 ();
 FILLCELL_X4 FILLER_144_557 ();
 FILLCELL_X1 FILLER_144_561 ();
 FILLCELL_X4 FILLER_144_584 ();
 FILLCELL_X1 FILLER_144_588 ();
 FILLCELL_X4 FILLER_144_596 ();
 FILLCELL_X2 FILLER_144_600 ();
 FILLCELL_X16 FILLER_144_614 ();
 FILLCELL_X1 FILLER_144_630 ();
 FILLCELL_X32 FILLER_144_632 ();
 FILLCELL_X16 FILLER_144_664 ();
 FILLCELL_X4 FILLER_144_680 ();
 FILLCELL_X1 FILLER_144_684 ();
 FILLCELL_X2 FILLER_144_705 ();
 FILLCELL_X4 FILLER_144_717 ();
 FILLCELL_X2 FILLER_144_721 ();
 FILLCELL_X2 FILLER_144_735 ();
 FILLCELL_X4 FILLER_144_755 ();
 FILLCELL_X2 FILLER_144_769 ();
 FILLCELL_X8 FILLER_144_782 ();
 FILLCELL_X4 FILLER_144_790 ();
 FILLCELL_X2 FILLER_144_794 ();
 FILLCELL_X8 FILLER_144_811 ();
 FILLCELL_X1 FILLER_144_819 ();
 FILLCELL_X2 FILLER_144_828 ();
 FILLCELL_X1 FILLER_144_834 ();
 FILLCELL_X2 FILLER_144_846 ();
 FILLCELL_X8 FILLER_144_862 ();
 FILLCELL_X32 FILLER_144_885 ();
 FILLCELL_X4 FILLER_144_917 ();
 FILLCELL_X1 FILLER_144_921 ();
 FILLCELL_X4 FILLER_144_929 ();
 FILLCELL_X2 FILLER_144_933 ();
 FILLCELL_X1 FILLER_144_935 ();
 FILLCELL_X16 FILLER_144_953 ();
 FILLCELL_X2 FILLER_144_969 ();
 FILLCELL_X4 FILLER_144_1028 ();
 FILLCELL_X4 FILLER_144_1038 ();
 FILLCELL_X2 FILLER_144_1042 ();
 FILLCELL_X1 FILLER_144_1044 ();
 FILLCELL_X2 FILLER_144_1049 ();
 FILLCELL_X8 FILLER_144_1056 ();
 FILLCELL_X4 FILLER_144_1064 ();
 FILLCELL_X2 FILLER_144_1068 ();
 FILLCELL_X1 FILLER_144_1070 ();
 FILLCELL_X2 FILLER_144_1075 ();
 FILLCELL_X16 FILLER_144_1080 ();
 FILLCELL_X1 FILLER_144_1096 ();
 FILLCELL_X2 FILLER_144_1111 ();
 FILLCELL_X2 FILLER_144_1117 ();
 FILLCELL_X1 FILLER_144_1130 ();
 FILLCELL_X32 FILLER_144_1135 ();
 FILLCELL_X32 FILLER_144_1167 ();
 FILLCELL_X8 FILLER_144_1199 ();
 FILLCELL_X2 FILLER_144_1207 ();
 FILLCELL_X32 FILLER_145_1 ();
 FILLCELL_X32 FILLER_145_33 ();
 FILLCELL_X32 FILLER_145_65 ();
 FILLCELL_X32 FILLER_145_97 ();
 FILLCELL_X32 FILLER_145_129 ();
 FILLCELL_X32 FILLER_145_161 ();
 FILLCELL_X16 FILLER_145_193 ();
 FILLCELL_X2 FILLER_145_209 ();
 FILLCELL_X2 FILLER_145_233 ();
 FILLCELL_X2 FILLER_145_245 ();
 FILLCELL_X1 FILLER_145_254 ();
 FILLCELL_X1 FILLER_145_261 ();
 FILLCELL_X4 FILLER_145_269 ();
 FILLCELL_X1 FILLER_145_273 ();
 FILLCELL_X16 FILLER_145_305 ();
 FILLCELL_X4 FILLER_145_321 ();
 FILLCELL_X1 FILLER_145_325 ();
 FILLCELL_X8 FILLER_145_330 ();
 FILLCELL_X1 FILLER_145_345 ();
 FILLCELL_X16 FILLER_145_350 ();
 FILLCELL_X2 FILLER_145_369 ();
 FILLCELL_X4 FILLER_145_380 ();
 FILLCELL_X1 FILLER_145_384 ();
 FILLCELL_X32 FILLER_145_390 ();
 FILLCELL_X16 FILLER_145_422 ();
 FILLCELL_X1 FILLER_145_438 ();
 FILLCELL_X1 FILLER_145_454 ();
 FILLCELL_X8 FILLER_145_477 ();
 FILLCELL_X1 FILLER_145_485 ();
 FILLCELL_X1 FILLER_145_505 ();
 FILLCELL_X8 FILLER_145_517 ();
 FILLCELL_X2 FILLER_145_525 ();
 FILLCELL_X1 FILLER_145_558 ();
 FILLCELL_X2 FILLER_145_564 ();
 FILLCELL_X1 FILLER_145_566 ();
 FILLCELL_X32 FILLER_145_631 ();
 FILLCELL_X16 FILLER_145_663 ();
 FILLCELL_X4 FILLER_145_679 ();
 FILLCELL_X2 FILLER_145_683 ();
 FILLCELL_X4 FILLER_145_692 ();
 FILLCELL_X2 FILLER_145_707 ();
 FILLCELL_X1 FILLER_145_724 ();
 FILLCELL_X4 FILLER_145_732 ();
 FILLCELL_X2 FILLER_145_736 ();
 FILLCELL_X1 FILLER_145_741 ();
 FILLCELL_X1 FILLER_145_757 ();
 FILLCELL_X8 FILLER_145_766 ();
 FILLCELL_X4 FILLER_145_774 ();
 FILLCELL_X2 FILLER_145_778 ();
 FILLCELL_X1 FILLER_145_780 ();
 FILLCELL_X1 FILLER_145_795 ();
 FILLCELL_X2 FILLER_145_807 ();
 FILLCELL_X2 FILLER_145_835 ();
 FILLCELL_X1 FILLER_145_871 ();
 FILLCELL_X2 FILLER_145_875 ();
 FILLCELL_X1 FILLER_145_877 ();
 FILLCELL_X32 FILLER_145_882 ();
 FILLCELL_X32 FILLER_145_914 ();
 FILLCELL_X16 FILLER_145_946 ();
 FILLCELL_X2 FILLER_145_962 ();
 FILLCELL_X1 FILLER_145_964 ();
 FILLCELL_X1 FILLER_145_976 ();
 FILLCELL_X2 FILLER_145_984 ();
 FILLCELL_X2 FILLER_145_1004 ();
 FILLCELL_X1 FILLER_145_1006 ();
 FILLCELL_X8 FILLER_145_1011 ();
 FILLCELL_X8 FILLER_145_1028 ();
 FILLCELL_X2 FILLER_145_1036 ();
 FILLCELL_X1 FILLER_145_1038 ();
 FILLCELL_X2 FILLER_145_1057 ();
 FILLCELL_X8 FILLER_145_1074 ();
 FILLCELL_X2 FILLER_145_1095 ();
 FILLCELL_X1 FILLER_145_1097 ();
 FILLCELL_X2 FILLER_145_1110 ();
 FILLCELL_X1 FILLER_145_1112 ();
 FILLCELL_X2 FILLER_145_1118 ();
 FILLCELL_X2 FILLER_145_1124 ();
 FILLCELL_X1 FILLER_145_1126 ();
 FILLCELL_X32 FILLER_145_1131 ();
 FILLCELL_X32 FILLER_145_1163 ();
 FILLCELL_X8 FILLER_145_1195 ();
 FILLCELL_X4 FILLER_145_1203 ();
 FILLCELL_X2 FILLER_145_1207 ();
 FILLCELL_X32 FILLER_146_1 ();
 FILLCELL_X32 FILLER_146_33 ();
 FILLCELL_X32 FILLER_146_65 ();
 FILLCELL_X32 FILLER_146_97 ();
 FILLCELL_X32 FILLER_146_129 ();
 FILLCELL_X32 FILLER_146_161 ();
 FILLCELL_X16 FILLER_146_193 ();
 FILLCELL_X4 FILLER_146_209 ();
 FILLCELL_X1 FILLER_146_213 ();
 FILLCELL_X2 FILLER_146_224 ();
 FILLCELL_X2 FILLER_146_269 ();
 FILLCELL_X2 FILLER_146_284 ();
 FILLCELL_X1 FILLER_146_286 ();
 FILLCELL_X4 FILLER_146_317 ();
 FILLCELL_X2 FILLER_146_321 ();
 FILLCELL_X1 FILLER_146_327 ();
 FILLCELL_X1 FILLER_146_335 ();
 FILLCELL_X2 FILLER_146_340 ();
 FILLCELL_X2 FILLER_146_345 ();
 FILLCELL_X1 FILLER_146_347 ();
 FILLCELL_X2 FILLER_146_372 ();
 FILLCELL_X2 FILLER_146_378 ();
 FILLCELL_X1 FILLER_146_380 ();
 FILLCELL_X2 FILLER_146_390 ();
 FILLCELL_X32 FILLER_146_398 ();
 FILLCELL_X2 FILLER_146_430 ();
 FILLCELL_X1 FILLER_146_432 ();
 FILLCELL_X4 FILLER_146_461 ();
 FILLCELL_X1 FILLER_146_469 ();
 FILLCELL_X2 FILLER_146_477 ();
 FILLCELL_X1 FILLER_146_479 ();
 FILLCELL_X8 FILLER_146_484 ();
 FILLCELL_X1 FILLER_146_492 ();
 FILLCELL_X4 FILLER_146_497 ();
 FILLCELL_X2 FILLER_146_501 ();
 FILLCELL_X2 FILLER_146_507 ();
 FILLCELL_X2 FILLER_146_517 ();
 FILLCELL_X1 FILLER_146_519 ();
 FILLCELL_X1 FILLER_146_524 ();
 FILLCELL_X1 FILLER_146_529 ();
 FILLCELL_X1 FILLER_146_545 ();
 FILLCELL_X1 FILLER_146_557 ();
 FILLCELL_X1 FILLER_146_562 ();
 FILLCELL_X8 FILLER_146_616 ();
 FILLCELL_X4 FILLER_146_624 ();
 FILLCELL_X2 FILLER_146_628 ();
 FILLCELL_X1 FILLER_146_630 ();
 FILLCELL_X32 FILLER_146_632 ();
 FILLCELL_X16 FILLER_146_664 ();
 FILLCELL_X2 FILLER_146_680 ();
 FILLCELL_X1 FILLER_146_682 ();
 FILLCELL_X4 FILLER_146_697 ();
 FILLCELL_X2 FILLER_146_701 ();
 FILLCELL_X4 FILLER_146_708 ();
 FILLCELL_X8 FILLER_146_736 ();
 FILLCELL_X4 FILLER_146_744 ();
 FILLCELL_X2 FILLER_146_748 ();
 FILLCELL_X4 FILLER_146_754 ();
 FILLCELL_X8 FILLER_146_773 ();
 FILLCELL_X4 FILLER_146_781 ();
 FILLCELL_X1 FILLER_146_789 ();
 FILLCELL_X8 FILLER_146_793 ();
 FILLCELL_X4 FILLER_146_801 ();
 FILLCELL_X1 FILLER_146_805 ();
 FILLCELL_X2 FILLER_146_812 ();
 FILLCELL_X1 FILLER_146_814 ();
 FILLCELL_X2 FILLER_146_847 ();
 FILLCELL_X1 FILLER_146_849 ();
 FILLCELL_X2 FILLER_146_865 ();
 FILLCELL_X1 FILLER_146_867 ();
 FILLCELL_X32 FILLER_146_891 ();
 FILLCELL_X32 FILLER_146_923 ();
 FILLCELL_X1 FILLER_146_955 ();
 FILLCELL_X1 FILLER_146_985 ();
 FILLCELL_X1 FILLER_146_1012 ();
 FILLCELL_X2 FILLER_146_1017 ();
 FILLCELL_X1 FILLER_146_1022 ();
 FILLCELL_X1 FILLER_146_1034 ();
 FILLCELL_X16 FILLER_146_1044 ();
 FILLCELL_X8 FILLER_146_1060 ();
 FILLCELL_X2 FILLER_146_1068 ();
 FILLCELL_X1 FILLER_146_1075 ();
 FILLCELL_X2 FILLER_146_1079 ();
 FILLCELL_X8 FILLER_146_1084 ();
 FILLCELL_X4 FILLER_146_1092 ();
 FILLCELL_X1 FILLER_146_1096 ();
 FILLCELL_X4 FILLER_146_1101 ();
 FILLCELL_X1 FILLER_146_1105 ();
 FILLCELL_X32 FILLER_146_1124 ();
 FILLCELL_X32 FILLER_146_1156 ();
 FILLCELL_X16 FILLER_146_1188 ();
 FILLCELL_X4 FILLER_146_1204 ();
 FILLCELL_X1 FILLER_146_1208 ();
 FILLCELL_X32 FILLER_147_1 ();
 FILLCELL_X32 FILLER_147_33 ();
 FILLCELL_X32 FILLER_147_65 ();
 FILLCELL_X32 FILLER_147_97 ();
 FILLCELL_X32 FILLER_147_129 ();
 FILLCELL_X32 FILLER_147_161 ();
 FILLCELL_X32 FILLER_147_193 ();
 FILLCELL_X1 FILLER_147_252 ();
 FILLCELL_X1 FILLER_147_262 ();
 FILLCELL_X2 FILLER_147_266 ();
 FILLCELL_X4 FILLER_147_273 ();
 FILLCELL_X2 FILLER_147_307 ();
 FILLCELL_X2 FILLER_147_317 ();
 FILLCELL_X2 FILLER_147_322 ();
 FILLCELL_X1 FILLER_147_324 ();
 FILLCELL_X4 FILLER_147_330 ();
 FILLCELL_X4 FILLER_147_344 ();
 FILLCELL_X2 FILLER_147_348 ();
 FILLCELL_X4 FILLER_147_355 ();
 FILLCELL_X2 FILLER_147_359 ();
 FILLCELL_X1 FILLER_147_361 ();
 FILLCELL_X1 FILLER_147_368 ();
 FILLCELL_X32 FILLER_147_399 ();
 FILLCELL_X8 FILLER_147_431 ();
 FILLCELL_X4 FILLER_147_439 ();
 FILLCELL_X2 FILLER_147_443 ();
 FILLCELL_X2 FILLER_147_449 ();
 FILLCELL_X1 FILLER_147_451 ();
 FILLCELL_X4 FILLER_147_456 ();
 FILLCELL_X2 FILLER_147_460 ();
 FILLCELL_X1 FILLER_147_462 ();
 FILLCELL_X1 FILLER_147_479 ();
 FILLCELL_X4 FILLER_147_484 ();
 FILLCELL_X2 FILLER_147_488 ();
 FILLCELL_X1 FILLER_147_490 ();
 FILLCELL_X2 FILLER_147_495 ();
 FILLCELL_X4 FILLER_147_501 ();
 FILLCELL_X2 FILLER_147_505 ();
 FILLCELL_X1 FILLER_147_507 ();
 FILLCELL_X16 FILLER_147_516 ();
 FILLCELL_X2 FILLER_147_532 ();
 FILLCELL_X1 FILLER_147_534 ();
 FILLCELL_X2 FILLER_147_542 ();
 FILLCELL_X2 FILLER_147_547 ();
 FILLCELL_X1 FILLER_147_556 ();
 FILLCELL_X2 FILLER_147_588 ();
 FILLCELL_X32 FILLER_147_626 ();
 FILLCELL_X8 FILLER_147_658 ();
 FILLCELL_X4 FILLER_147_666 ();
 FILLCELL_X2 FILLER_147_670 ();
 FILLCELL_X1 FILLER_147_672 ();
 FILLCELL_X4 FILLER_147_695 ();
 FILLCELL_X1 FILLER_147_699 ();
 FILLCELL_X2 FILLER_147_704 ();
 FILLCELL_X1 FILLER_147_706 ();
 FILLCELL_X4 FILLER_147_721 ();
 FILLCELL_X4 FILLER_147_729 ();
 FILLCELL_X2 FILLER_147_733 ();
 FILLCELL_X2 FILLER_147_780 ();
 FILLCELL_X2 FILLER_147_794 ();
 FILLCELL_X4 FILLER_147_811 ();
 FILLCELL_X2 FILLER_147_815 ();
 FILLCELL_X1 FILLER_147_817 ();
 FILLCELL_X32 FILLER_147_888 ();
 FILLCELL_X32 FILLER_147_920 ();
 FILLCELL_X16 FILLER_147_952 ();
 FILLCELL_X8 FILLER_147_968 ();
 FILLCELL_X2 FILLER_147_976 ();
 FILLCELL_X1 FILLER_147_978 ();
 FILLCELL_X2 FILLER_147_986 ();
 FILLCELL_X1 FILLER_147_988 ();
 FILLCELL_X8 FILLER_147_993 ();
 FILLCELL_X4 FILLER_147_1001 ();
 FILLCELL_X8 FILLER_147_1012 ();
 FILLCELL_X4 FILLER_147_1020 ();
 FILLCELL_X2 FILLER_147_1024 ();
 FILLCELL_X1 FILLER_147_1026 ();
 FILLCELL_X2 FILLER_147_1055 ();
 FILLCELL_X1 FILLER_147_1057 ();
 FILLCELL_X1 FILLER_147_1061 ();
 FILLCELL_X2 FILLER_147_1069 ();
 FILLCELL_X8 FILLER_147_1086 ();
 FILLCELL_X8 FILLER_147_1098 ();
 FILLCELL_X1 FILLER_147_1121 ();
 FILLCELL_X32 FILLER_147_1129 ();
 FILLCELL_X32 FILLER_147_1161 ();
 FILLCELL_X16 FILLER_147_1193 ();
 FILLCELL_X32 FILLER_148_1 ();
 FILLCELL_X32 FILLER_148_33 ();
 FILLCELL_X32 FILLER_148_65 ();
 FILLCELL_X32 FILLER_148_97 ();
 FILLCELL_X32 FILLER_148_129 ();
 FILLCELL_X32 FILLER_148_161 ();
 FILLCELL_X16 FILLER_148_193 ();
 FILLCELL_X4 FILLER_148_219 ();
 FILLCELL_X2 FILLER_148_223 ();
 FILLCELL_X1 FILLER_148_225 ();
 FILLCELL_X1 FILLER_148_233 ();
 FILLCELL_X1 FILLER_148_241 ();
 FILLCELL_X2 FILLER_148_249 ();
 FILLCELL_X1 FILLER_148_251 ();
 FILLCELL_X2 FILLER_148_260 ();
 FILLCELL_X8 FILLER_148_270 ();
 FILLCELL_X2 FILLER_148_278 ();
 FILLCELL_X4 FILLER_148_283 ();
 FILLCELL_X2 FILLER_148_287 ();
 FILLCELL_X1 FILLER_148_289 ();
 FILLCELL_X8 FILLER_148_300 ();
 FILLCELL_X1 FILLER_148_308 ();
 FILLCELL_X2 FILLER_148_329 ();
 FILLCELL_X1 FILLER_148_331 ();
 FILLCELL_X2 FILLER_148_347 ();
 FILLCELL_X1 FILLER_148_349 ();
 FILLCELL_X2 FILLER_148_358 ();
 FILLCELL_X1 FILLER_148_360 ();
 FILLCELL_X2 FILLER_148_365 ();
 FILLCELL_X1 FILLER_148_384 ();
 FILLCELL_X1 FILLER_148_389 ();
 FILLCELL_X32 FILLER_148_397 ();
 FILLCELL_X16 FILLER_148_429 ();
 FILLCELL_X4 FILLER_148_445 ();
 FILLCELL_X2 FILLER_148_460 ();
 FILLCELL_X1 FILLER_148_462 ();
 FILLCELL_X1 FILLER_148_470 ();
 FILLCELL_X1 FILLER_148_496 ();
 FILLCELL_X4 FILLER_148_507 ();
 FILLCELL_X4 FILLER_148_525 ();
 FILLCELL_X4 FILLER_148_536 ();
 FILLCELL_X2 FILLER_148_563 ();
 FILLCELL_X8 FILLER_148_569 ();
 FILLCELL_X2 FILLER_148_577 ();
 FILLCELL_X1 FILLER_148_592 ();
 FILLCELL_X16 FILLER_148_605 ();
 FILLCELL_X8 FILLER_148_621 ();
 FILLCELL_X2 FILLER_148_629 ();
 FILLCELL_X32 FILLER_148_632 ();
 FILLCELL_X16 FILLER_148_664 ();
 FILLCELL_X4 FILLER_148_680 ();
 FILLCELL_X2 FILLER_148_684 ();
 FILLCELL_X4 FILLER_148_700 ();
 FILLCELL_X2 FILLER_148_744 ();
 FILLCELL_X2 FILLER_148_756 ();
 FILLCELL_X1 FILLER_148_771 ();
 FILLCELL_X1 FILLER_148_784 ();
 FILLCELL_X16 FILLER_148_791 ();
 FILLCELL_X2 FILLER_148_807 ();
 FILLCELL_X1 FILLER_148_809 ();
 FILLCELL_X4 FILLER_148_831 ();
 FILLCELL_X2 FILLER_148_842 ();
 FILLCELL_X1 FILLER_148_844 ();
 FILLCELL_X1 FILLER_148_873 ();
 FILLCELL_X32 FILLER_148_886 ();
 FILLCELL_X32 FILLER_148_918 ();
 FILLCELL_X2 FILLER_148_950 ();
 FILLCELL_X8 FILLER_148_965 ();
 FILLCELL_X2 FILLER_148_973 ();
 FILLCELL_X1 FILLER_148_975 ();
 FILLCELL_X2 FILLER_148_1002 ();
 FILLCELL_X2 FILLER_148_1025 ();
 FILLCELL_X1 FILLER_148_1048 ();
 FILLCELL_X1 FILLER_148_1053 ();
 FILLCELL_X2 FILLER_148_1059 ();
 FILLCELL_X4 FILLER_148_1072 ();
 FILLCELL_X2 FILLER_148_1076 ();
 FILLCELL_X1 FILLER_148_1078 ();
 FILLCELL_X2 FILLER_148_1105 ();
 FILLCELL_X2 FILLER_148_1116 ();
 FILLCELL_X1 FILLER_148_1118 ();
 FILLCELL_X4 FILLER_148_1123 ();
 FILLCELL_X32 FILLER_148_1138 ();
 FILLCELL_X32 FILLER_148_1170 ();
 FILLCELL_X4 FILLER_148_1202 ();
 FILLCELL_X2 FILLER_148_1206 ();
 FILLCELL_X1 FILLER_148_1208 ();
 FILLCELL_X32 FILLER_149_1 ();
 FILLCELL_X32 FILLER_149_33 ();
 FILLCELL_X32 FILLER_149_65 ();
 FILLCELL_X32 FILLER_149_97 ();
 FILLCELL_X32 FILLER_149_129 ();
 FILLCELL_X32 FILLER_149_161 ();
 FILLCELL_X16 FILLER_149_193 ();
 FILLCELL_X4 FILLER_149_209 ();
 FILLCELL_X2 FILLER_149_213 ();
 FILLCELL_X2 FILLER_149_232 ();
 FILLCELL_X1 FILLER_149_234 ();
 FILLCELL_X2 FILLER_149_257 ();
 FILLCELL_X1 FILLER_149_259 ();
 FILLCELL_X1 FILLER_149_264 ();
 FILLCELL_X1 FILLER_149_272 ();
 FILLCELL_X2 FILLER_149_278 ();
 FILLCELL_X1 FILLER_149_287 ();
 FILLCELL_X4 FILLER_149_292 ();
 FILLCELL_X1 FILLER_149_296 ();
 FILLCELL_X4 FILLER_149_315 ();
 FILLCELL_X2 FILLER_149_319 ();
 FILLCELL_X2 FILLER_149_331 ();
 FILLCELL_X1 FILLER_149_333 ();
 FILLCELL_X1 FILLER_149_338 ();
 FILLCELL_X1 FILLER_149_345 ();
 FILLCELL_X2 FILLER_149_353 ();
 FILLCELL_X1 FILLER_149_362 ();
 FILLCELL_X2 FILLER_149_383 ();
 FILLCELL_X1 FILLER_149_385 ();
 FILLCELL_X32 FILLER_149_398 ();
 FILLCELL_X8 FILLER_149_430 ();
 FILLCELL_X4 FILLER_149_448 ();
 FILLCELL_X1 FILLER_149_452 ();
 FILLCELL_X2 FILLER_149_462 ();
 FILLCELL_X4 FILLER_149_468 ();
 FILLCELL_X1 FILLER_149_472 ();
 FILLCELL_X2 FILLER_149_494 ();
 FILLCELL_X1 FILLER_149_496 ();
 FILLCELL_X16 FILLER_149_519 ();
 FILLCELL_X1 FILLER_149_535 ();
 FILLCELL_X8 FILLER_149_547 ();
 FILLCELL_X2 FILLER_149_558 ();
 FILLCELL_X2 FILLER_149_567 ();
 FILLCELL_X1 FILLER_149_569 ();
 FILLCELL_X32 FILLER_149_617 ();
 FILLCELL_X32 FILLER_149_649 ();
 FILLCELL_X1 FILLER_149_681 ();
 FILLCELL_X2 FILLER_149_703 ();
 FILLCELL_X1 FILLER_149_705 ();
 FILLCELL_X1 FILLER_149_715 ();
 FILLCELL_X8 FILLER_149_732 ();
 FILLCELL_X1 FILLER_149_740 ();
 FILLCELL_X1 FILLER_149_745 ();
 FILLCELL_X1 FILLER_149_750 ();
 FILLCELL_X8 FILLER_149_755 ();
 FILLCELL_X4 FILLER_149_763 ();
 FILLCELL_X8 FILLER_149_770 ();
 FILLCELL_X4 FILLER_149_778 ();
 FILLCELL_X2 FILLER_149_782 ();
 FILLCELL_X1 FILLER_149_799 ();
 FILLCELL_X2 FILLER_149_804 ();
 FILLCELL_X4 FILLER_149_814 ();
 FILLCELL_X1 FILLER_149_821 ();
 FILLCELL_X8 FILLER_149_825 ();
 FILLCELL_X4 FILLER_149_833 ();
 FILLCELL_X1 FILLER_149_837 ();
 FILLCELL_X2 FILLER_149_849 ();
 FILLCELL_X1 FILLER_149_851 ();
 FILLCELL_X1 FILLER_149_860 ();
 FILLCELL_X1 FILLER_149_866 ();
 FILLCELL_X32 FILLER_149_876 ();
 FILLCELL_X32 FILLER_149_908 ();
 FILLCELL_X8 FILLER_149_940 ();
 FILLCELL_X4 FILLER_149_948 ();
 FILLCELL_X2 FILLER_149_952 ();
 FILLCELL_X1 FILLER_149_954 ();
 FILLCELL_X2 FILLER_149_968 ();
 FILLCELL_X2 FILLER_149_999 ();
 FILLCELL_X16 FILLER_149_1015 ();
 FILLCELL_X2 FILLER_149_1036 ();
 FILLCELL_X2 FILLER_149_1043 ();
 FILLCELL_X1 FILLER_149_1045 ();
 FILLCELL_X4 FILLER_149_1058 ();
 FILLCELL_X4 FILLER_149_1068 ();
 FILLCELL_X2 FILLER_149_1072 ();
 FILLCELL_X8 FILLER_149_1090 ();
 FILLCELL_X4 FILLER_149_1098 ();
 FILLCELL_X2 FILLER_149_1113 ();
 FILLCELL_X2 FILLER_149_1119 ();
 FILLCELL_X1 FILLER_149_1132 ();
 FILLCELL_X32 FILLER_149_1136 ();
 FILLCELL_X32 FILLER_149_1168 ();
 FILLCELL_X8 FILLER_149_1200 ();
 FILLCELL_X1 FILLER_149_1208 ();
 FILLCELL_X32 FILLER_150_1 ();
 FILLCELL_X32 FILLER_150_33 ();
 FILLCELL_X32 FILLER_150_65 ();
 FILLCELL_X32 FILLER_150_97 ();
 FILLCELL_X32 FILLER_150_129 ();
 FILLCELL_X32 FILLER_150_161 ();
 FILLCELL_X16 FILLER_150_193 ();
 FILLCELL_X4 FILLER_150_209 ();
 FILLCELL_X4 FILLER_150_230 ();
 FILLCELL_X1 FILLER_150_239 ();
 FILLCELL_X2 FILLER_150_244 ();
 FILLCELL_X8 FILLER_150_250 ();
 FILLCELL_X4 FILLER_150_258 ();
 FILLCELL_X2 FILLER_150_262 ();
 FILLCELL_X1 FILLER_150_264 ();
 FILLCELL_X1 FILLER_150_277 ();
 FILLCELL_X2 FILLER_150_293 ();
 FILLCELL_X1 FILLER_150_295 ();
 FILLCELL_X1 FILLER_150_305 ();
 FILLCELL_X1 FILLER_150_314 ();
 FILLCELL_X1 FILLER_150_341 ();
 FILLCELL_X1 FILLER_150_347 ();
 FILLCELL_X2 FILLER_150_354 ();
 FILLCELL_X4 FILLER_150_366 ();
 FILLCELL_X32 FILLER_150_395 ();
 FILLCELL_X8 FILLER_150_427 ();
 FILLCELL_X2 FILLER_150_435 ();
 FILLCELL_X1 FILLER_150_437 ();
 FILLCELL_X1 FILLER_150_457 ();
 FILLCELL_X2 FILLER_150_473 ();
 FILLCELL_X1 FILLER_150_475 ();
 FILLCELL_X8 FILLER_150_480 ();
 FILLCELL_X4 FILLER_150_488 ();
 FILLCELL_X2 FILLER_150_492 ();
 FILLCELL_X1 FILLER_150_494 ();
 FILLCELL_X4 FILLER_150_502 ();
 FILLCELL_X2 FILLER_150_506 ();
 FILLCELL_X1 FILLER_150_508 ();
 FILLCELL_X1 FILLER_150_522 ();
 FILLCELL_X1 FILLER_150_527 ();
 FILLCELL_X2 FILLER_150_532 ();
 FILLCELL_X1 FILLER_150_534 ();
 FILLCELL_X8 FILLER_150_546 ();
 FILLCELL_X1 FILLER_150_554 ();
 FILLCELL_X8 FILLER_150_569 ();
 FILLCELL_X1 FILLER_150_577 ();
 FILLCELL_X2 FILLER_150_597 ();
 FILLCELL_X1 FILLER_150_609 ();
 FILLCELL_X8 FILLER_150_617 ();
 FILLCELL_X4 FILLER_150_625 ();
 FILLCELL_X2 FILLER_150_629 ();
 FILLCELL_X32 FILLER_150_632 ();
 FILLCELL_X16 FILLER_150_664 ();
 FILLCELL_X8 FILLER_150_680 ();
 FILLCELL_X4 FILLER_150_688 ();
 FILLCELL_X4 FILLER_150_708 ();
 FILLCELL_X4 FILLER_150_729 ();
 FILLCELL_X4 FILLER_150_755 ();
 FILLCELL_X2 FILLER_150_763 ();
 FILLCELL_X4 FILLER_150_777 ();
 FILLCELL_X1 FILLER_150_781 ();
 FILLCELL_X4 FILLER_150_790 ();
 FILLCELL_X2 FILLER_150_794 ();
 FILLCELL_X1 FILLER_150_805 ();
 FILLCELL_X4 FILLER_150_823 ();
 FILLCELL_X1 FILLER_150_827 ();
 FILLCELL_X1 FILLER_150_834 ();
 FILLCELL_X2 FILLER_150_841 ();
 FILLCELL_X2 FILLER_150_851 ();
 FILLCELL_X1 FILLER_150_860 ();
 FILLCELL_X1 FILLER_150_864 ();
 FILLCELL_X1 FILLER_150_870 ();
 FILLCELL_X32 FILLER_150_875 ();
 FILLCELL_X32 FILLER_150_907 ();
 FILLCELL_X32 FILLER_150_939 ();
 FILLCELL_X16 FILLER_150_971 ();
 FILLCELL_X1 FILLER_150_987 ();
 FILLCELL_X4 FILLER_150_1002 ();
 FILLCELL_X8 FILLER_150_1062 ();
 FILLCELL_X8 FILLER_150_1090 ();
 FILLCELL_X4 FILLER_150_1112 ();
 FILLCELL_X2 FILLER_150_1116 ();
 FILLCELL_X2 FILLER_150_1127 ();
 FILLCELL_X1 FILLER_150_1129 ();
 FILLCELL_X32 FILLER_150_1139 ();
 FILLCELL_X32 FILLER_150_1171 ();
 FILLCELL_X4 FILLER_150_1203 ();
 FILLCELL_X2 FILLER_150_1207 ();
 FILLCELL_X32 FILLER_151_1 ();
 FILLCELL_X32 FILLER_151_33 ();
 FILLCELL_X32 FILLER_151_65 ();
 FILLCELL_X32 FILLER_151_97 ();
 FILLCELL_X32 FILLER_151_129 ();
 FILLCELL_X32 FILLER_151_161 ();
 FILLCELL_X32 FILLER_151_193 ();
 FILLCELL_X1 FILLER_151_225 ();
 FILLCELL_X2 FILLER_151_230 ();
 FILLCELL_X1 FILLER_151_232 ();
 FILLCELL_X2 FILLER_151_251 ();
 FILLCELL_X1 FILLER_151_253 ();
 FILLCELL_X4 FILLER_151_262 ();
 FILLCELL_X2 FILLER_151_266 ();
 FILLCELL_X8 FILLER_151_285 ();
 FILLCELL_X4 FILLER_151_293 ();
 FILLCELL_X1 FILLER_151_297 ();
 FILLCELL_X4 FILLER_151_306 ();
 FILLCELL_X1 FILLER_151_319 ();
 FILLCELL_X1 FILLER_151_326 ();
 FILLCELL_X2 FILLER_151_334 ();
 FILLCELL_X1 FILLER_151_340 ();
 FILLCELL_X1 FILLER_151_364 ();
 FILLCELL_X1 FILLER_151_368 ();
 FILLCELL_X1 FILLER_151_376 ();
 FILLCELL_X1 FILLER_151_381 ();
 FILLCELL_X32 FILLER_151_400 ();
 FILLCELL_X8 FILLER_151_432 ();
 FILLCELL_X1 FILLER_151_440 ();
 FILLCELL_X2 FILLER_151_462 ();
 FILLCELL_X2 FILLER_151_468 ();
 FILLCELL_X1 FILLER_151_470 ();
 FILLCELL_X2 FILLER_151_475 ();
 FILLCELL_X1 FILLER_151_477 ();
 FILLCELL_X2 FILLER_151_482 ();
 FILLCELL_X4 FILLER_151_498 ();
 FILLCELL_X2 FILLER_151_507 ();
 FILLCELL_X2 FILLER_151_518 ();
 FILLCELL_X16 FILLER_151_524 ();
 FILLCELL_X2 FILLER_151_540 ();
 FILLCELL_X1 FILLER_151_542 ();
 FILLCELL_X8 FILLER_151_546 ();
 FILLCELL_X2 FILLER_151_554 ();
 FILLCELL_X1 FILLER_151_556 ();
 FILLCELL_X4 FILLER_151_567 ();
 FILLCELL_X2 FILLER_151_571 ();
 FILLCELL_X1 FILLER_151_580 ();
 FILLCELL_X2 FILLER_151_601 ();
 FILLCELL_X1 FILLER_151_603 ();
 FILLCELL_X32 FILLER_151_627 ();
 FILLCELL_X16 FILLER_151_659 ();
 FILLCELL_X8 FILLER_151_675 ();
 FILLCELL_X1 FILLER_151_703 ();
 FILLCELL_X1 FILLER_151_730 ();
 FILLCELL_X1 FILLER_151_735 ();
 FILLCELL_X1 FILLER_151_743 ();
 FILLCELL_X8 FILLER_151_755 ();
 FILLCELL_X4 FILLER_151_763 ();
 FILLCELL_X4 FILLER_151_777 ();
 FILLCELL_X4 FILLER_151_789 ();
 FILLCELL_X1 FILLER_151_793 ();
 FILLCELL_X1 FILLER_151_798 ();
 FILLCELL_X8 FILLER_151_837 ();
 FILLCELL_X2 FILLER_151_856 ();
 FILLCELL_X4 FILLER_151_862 ();
 FILLCELL_X32 FILLER_151_880 ();
 FILLCELL_X32 FILLER_151_912 ();
 FILLCELL_X32 FILLER_151_944 ();
 FILLCELL_X4 FILLER_151_976 ();
 FILLCELL_X2 FILLER_151_980 ();
 FILLCELL_X1 FILLER_151_982 ();
 FILLCELL_X4 FILLER_151_990 ();
 FILLCELL_X2 FILLER_151_994 ();
 FILLCELL_X1 FILLER_151_1008 ();
 FILLCELL_X1 FILLER_151_1016 ();
 FILLCELL_X4 FILLER_151_1021 ();
 FILLCELL_X1 FILLER_151_1025 ();
 FILLCELL_X4 FILLER_151_1029 ();
 FILLCELL_X2 FILLER_151_1033 ();
 FILLCELL_X1 FILLER_151_1035 ();
 FILLCELL_X4 FILLER_151_1045 ();
 FILLCELL_X2 FILLER_151_1049 ();
 FILLCELL_X2 FILLER_151_1055 ();
 FILLCELL_X1 FILLER_151_1057 ();
 FILLCELL_X8 FILLER_151_1062 ();
 FILLCELL_X4 FILLER_151_1070 ();
 FILLCELL_X2 FILLER_151_1093 ();
 FILLCELL_X2 FILLER_151_1099 ();
 FILLCELL_X1 FILLER_151_1119 ();
 FILLCELL_X32 FILLER_151_1127 ();
 FILLCELL_X32 FILLER_151_1159 ();
 FILLCELL_X16 FILLER_151_1191 ();
 FILLCELL_X2 FILLER_151_1207 ();
 FILLCELL_X32 FILLER_152_1 ();
 FILLCELL_X32 FILLER_152_33 ();
 FILLCELL_X32 FILLER_152_65 ();
 FILLCELL_X32 FILLER_152_97 ();
 FILLCELL_X32 FILLER_152_129 ();
 FILLCELL_X32 FILLER_152_161 ();
 FILLCELL_X4 FILLER_152_193 ();
 FILLCELL_X2 FILLER_152_197 ();
 FILLCELL_X1 FILLER_152_199 ();
 FILLCELL_X4 FILLER_152_210 ();
 FILLCELL_X1 FILLER_152_214 ();
 FILLCELL_X4 FILLER_152_222 ();
 FILLCELL_X1 FILLER_152_226 ();
 FILLCELL_X2 FILLER_152_231 ();
 FILLCELL_X4 FILLER_152_240 ();
 FILLCELL_X4 FILLER_152_248 ();
 FILLCELL_X2 FILLER_152_252 ();
 FILLCELL_X2 FILLER_152_258 ();
 FILLCELL_X4 FILLER_152_264 ();
 FILLCELL_X8 FILLER_152_271 ();
 FILLCELL_X2 FILLER_152_279 ();
 FILLCELL_X2 FILLER_152_296 ();
 FILLCELL_X1 FILLER_152_298 ();
 FILLCELL_X2 FILLER_152_302 ();
 FILLCELL_X2 FILLER_152_311 ();
 FILLCELL_X1 FILLER_152_317 ();
 FILLCELL_X4 FILLER_152_325 ();
 FILLCELL_X4 FILLER_152_340 ();
 FILLCELL_X1 FILLER_152_344 ();
 FILLCELL_X1 FILLER_152_381 ();
 FILLCELL_X1 FILLER_152_393 ();
 FILLCELL_X32 FILLER_152_403 ();
 FILLCELL_X4 FILLER_152_435 ();
 FILLCELL_X2 FILLER_152_439 ();
 FILLCELL_X1 FILLER_152_441 ();
 FILLCELL_X8 FILLER_152_500 ();
 FILLCELL_X1 FILLER_152_508 ();
 FILLCELL_X2 FILLER_152_516 ();
 FILLCELL_X1 FILLER_152_518 ();
 FILLCELL_X4 FILLER_152_523 ();
 FILLCELL_X2 FILLER_152_527 ();
 FILLCELL_X1 FILLER_152_529 ();
 FILLCELL_X2 FILLER_152_533 ();
 FILLCELL_X8 FILLER_152_540 ();
 FILLCELL_X4 FILLER_152_548 ();
 FILLCELL_X1 FILLER_152_560 ();
 FILLCELL_X2 FILLER_152_568 ();
 FILLCELL_X1 FILLER_152_570 ();
 FILLCELL_X8 FILLER_152_619 ();
 FILLCELL_X4 FILLER_152_627 ();
 FILLCELL_X32 FILLER_152_632 ();
 FILLCELL_X16 FILLER_152_664 ();
 FILLCELL_X2 FILLER_152_680 ();
 FILLCELL_X8 FILLER_152_709 ();
 FILLCELL_X1 FILLER_152_717 ();
 FILLCELL_X2 FILLER_152_725 ();
 FILLCELL_X1 FILLER_152_727 ();
 FILLCELL_X2 FILLER_152_733 ();
 FILLCELL_X2 FILLER_152_739 ();
 FILLCELL_X1 FILLER_152_757 ();
 FILLCELL_X4 FILLER_152_765 ();
 FILLCELL_X2 FILLER_152_769 ();
 FILLCELL_X4 FILLER_152_778 ();
 FILLCELL_X2 FILLER_152_782 ();
 FILLCELL_X1 FILLER_152_784 ();
 FILLCELL_X8 FILLER_152_796 ();
 FILLCELL_X2 FILLER_152_804 ();
 FILLCELL_X2 FILLER_152_815 ();
 FILLCELL_X4 FILLER_152_821 ();
 FILLCELL_X1 FILLER_152_825 ();
 FILLCELL_X1 FILLER_152_829 ();
 FILLCELL_X1 FILLER_152_837 ();
 FILLCELL_X2 FILLER_152_844 ();
 FILLCELL_X2 FILLER_152_850 ();
 FILLCELL_X4 FILLER_152_857 ();
 FILLCELL_X1 FILLER_152_865 ();
 FILLCELL_X32 FILLER_152_877 ();
 FILLCELL_X32 FILLER_152_909 ();
 FILLCELL_X32 FILLER_152_941 ();
 FILLCELL_X16 FILLER_152_973 ();
 FILLCELL_X4 FILLER_152_989 ();
 FILLCELL_X2 FILLER_152_993 ();
 FILLCELL_X2 FILLER_152_1034 ();
 FILLCELL_X1 FILLER_152_1073 ();
 FILLCELL_X1 FILLER_152_1096 ();
 FILLCELL_X4 FILLER_152_1104 ();
 FILLCELL_X2 FILLER_152_1108 ();
 FILLCELL_X1 FILLER_152_1110 ();
 FILLCELL_X32 FILLER_152_1160 ();
 FILLCELL_X16 FILLER_152_1192 ();
 FILLCELL_X1 FILLER_152_1208 ();
 FILLCELL_X32 FILLER_153_1 ();
 FILLCELL_X32 FILLER_153_33 ();
 FILLCELL_X32 FILLER_153_65 ();
 FILLCELL_X32 FILLER_153_97 ();
 FILLCELL_X32 FILLER_153_129 ();
 FILLCELL_X32 FILLER_153_161 ();
 FILLCELL_X16 FILLER_153_193 ();
 FILLCELL_X2 FILLER_153_209 ();
 FILLCELL_X4 FILLER_153_238 ();
 FILLCELL_X1 FILLER_153_242 ();
 FILLCELL_X8 FILLER_153_279 ();
 FILLCELL_X4 FILLER_153_287 ();
 FILLCELL_X1 FILLER_153_291 ();
 FILLCELL_X16 FILLER_153_308 ();
 FILLCELL_X1 FILLER_153_324 ();
 FILLCELL_X1 FILLER_153_331 ();
 FILLCELL_X4 FILLER_153_335 ();
 FILLCELL_X1 FILLER_153_339 ();
 FILLCELL_X2 FILLER_153_344 ();
 FILLCELL_X1 FILLER_153_357 ();
 FILLCELL_X1 FILLER_153_388 ();
 FILLCELL_X2 FILLER_153_394 ();
 FILLCELL_X32 FILLER_153_400 ();
 FILLCELL_X4 FILLER_153_432 ();
 FILLCELL_X1 FILLER_153_436 ();
 FILLCELL_X2 FILLER_153_466 ();
 FILLCELL_X1 FILLER_153_472 ();
 FILLCELL_X4 FILLER_153_483 ();
 FILLCELL_X8 FILLER_153_494 ();
 FILLCELL_X4 FILLER_153_502 ();
 FILLCELL_X2 FILLER_153_506 ();
 FILLCELL_X4 FILLER_153_529 ();
 FILLCELL_X2 FILLER_153_554 ();
 FILLCELL_X2 FILLER_153_566 ();
 FILLCELL_X1 FILLER_153_568 ();
 FILLCELL_X2 FILLER_153_590 ();
 FILLCELL_X1 FILLER_153_592 ();
 FILLCELL_X32 FILLER_153_622 ();
 FILLCELL_X32 FILLER_153_654 ();
 FILLCELL_X8 FILLER_153_686 ();
 FILLCELL_X4 FILLER_153_694 ();
 FILLCELL_X2 FILLER_153_698 ();
 FILLCELL_X1 FILLER_153_700 ();
 FILLCELL_X2 FILLER_153_733 ();
 FILLCELL_X2 FILLER_153_777 ();
 FILLCELL_X2 FILLER_153_798 ();
 FILLCELL_X1 FILLER_153_800 ();
 FILLCELL_X1 FILLER_153_808 ();
 FILLCELL_X1 FILLER_153_830 ();
 FILLCELL_X4 FILLER_153_841 ();
 FILLCELL_X4 FILLER_153_850 ();
 FILLCELL_X32 FILLER_153_876 ();
 FILLCELL_X32 FILLER_153_908 ();
 FILLCELL_X32 FILLER_153_940 ();
 FILLCELL_X32 FILLER_153_972 ();
 FILLCELL_X32 FILLER_153_1004 ();
 FILLCELL_X8 FILLER_153_1036 ();
 FILLCELL_X1 FILLER_153_1044 ();
 FILLCELL_X1 FILLER_153_1052 ();
 FILLCELL_X32 FILLER_153_1060 ();
 FILLCELL_X32 FILLER_153_1092 ();
 FILLCELL_X32 FILLER_153_1124 ();
 FILLCELL_X32 FILLER_153_1156 ();
 FILLCELL_X16 FILLER_153_1188 ();
 FILLCELL_X4 FILLER_153_1204 ();
 FILLCELL_X1 FILLER_153_1208 ();
 FILLCELL_X32 FILLER_154_1 ();
 FILLCELL_X32 FILLER_154_33 ();
 FILLCELL_X32 FILLER_154_65 ();
 FILLCELL_X32 FILLER_154_97 ();
 FILLCELL_X32 FILLER_154_129 ();
 FILLCELL_X32 FILLER_154_161 ();
 FILLCELL_X32 FILLER_154_193 ();
 FILLCELL_X2 FILLER_154_225 ();
 FILLCELL_X1 FILLER_154_227 ();
 FILLCELL_X1 FILLER_154_238 ();
 FILLCELL_X4 FILLER_154_246 ();
 FILLCELL_X1 FILLER_154_250 ();
 FILLCELL_X2 FILLER_154_262 ();
 FILLCELL_X4 FILLER_154_270 ();
 FILLCELL_X8 FILLER_154_287 ();
 FILLCELL_X1 FILLER_154_295 ();
 FILLCELL_X1 FILLER_154_300 ();
 FILLCELL_X1 FILLER_154_307 ();
 FILLCELL_X1 FILLER_154_312 ();
 FILLCELL_X1 FILLER_154_320 ();
 FILLCELL_X4 FILLER_154_329 ();
 FILLCELL_X2 FILLER_154_339 ();
 FILLCELL_X1 FILLER_154_341 ();
 FILLCELL_X1 FILLER_154_363 ();
 FILLCELL_X4 FILLER_154_385 ();
 FILLCELL_X32 FILLER_154_394 ();
 FILLCELL_X16 FILLER_154_426 ();
 FILLCELL_X8 FILLER_154_442 ();
 FILLCELL_X4 FILLER_154_450 ();
 FILLCELL_X1 FILLER_154_454 ();
 FILLCELL_X2 FILLER_154_458 ();
 FILLCELL_X1 FILLER_154_460 ();
 FILLCELL_X4 FILLER_154_466 ();
 FILLCELL_X1 FILLER_154_470 ();
 FILLCELL_X1 FILLER_154_500 ();
 FILLCELL_X2 FILLER_154_508 ();
 FILLCELL_X2 FILLER_154_545 ();
 FILLCELL_X1 FILLER_154_547 ();
 FILLCELL_X2 FILLER_154_561 ();
 FILLCELL_X1 FILLER_154_574 ();
 FILLCELL_X2 FILLER_154_598 ();
 FILLCELL_X16 FILLER_154_611 ();
 FILLCELL_X4 FILLER_154_627 ();
 FILLCELL_X32 FILLER_154_632 ();
 FILLCELL_X16 FILLER_154_664 ();
 FILLCELL_X2 FILLER_154_680 ();
 FILLCELL_X1 FILLER_154_682 ();
 FILLCELL_X2 FILLER_154_693 ();
 FILLCELL_X2 FILLER_154_702 ();
 FILLCELL_X1 FILLER_154_704 ();
 FILLCELL_X4 FILLER_154_715 ();
 FILLCELL_X2 FILLER_154_746 ();
 FILLCELL_X2 FILLER_154_756 ();
 FILLCELL_X16 FILLER_154_777 ();
 FILLCELL_X4 FILLER_154_793 ();
 FILLCELL_X1 FILLER_154_797 ();
 FILLCELL_X8 FILLER_154_809 ();
 FILLCELL_X4 FILLER_154_817 ();
 FILLCELL_X2 FILLER_154_821 ();
 FILLCELL_X1 FILLER_154_823 ();
 FILLCELL_X1 FILLER_154_832 ();
 FILLCELL_X2 FILLER_154_837 ();
 FILLCELL_X32 FILLER_154_875 ();
 FILLCELL_X32 FILLER_154_907 ();
 FILLCELL_X32 FILLER_154_939 ();
 FILLCELL_X32 FILLER_154_971 ();
 FILLCELL_X32 FILLER_154_1003 ();
 FILLCELL_X8 FILLER_154_1035 ();
 FILLCELL_X4 FILLER_154_1043 ();
 FILLCELL_X2 FILLER_154_1047 ();
 FILLCELL_X32 FILLER_154_1062 ();
 FILLCELL_X32 FILLER_154_1094 ();
 FILLCELL_X32 FILLER_154_1126 ();
 FILLCELL_X32 FILLER_154_1158 ();
 FILLCELL_X16 FILLER_154_1190 ();
 FILLCELL_X2 FILLER_154_1206 ();
 FILLCELL_X1 FILLER_154_1208 ();
 FILLCELL_X32 FILLER_155_1 ();
 FILLCELL_X32 FILLER_155_33 ();
 FILLCELL_X32 FILLER_155_65 ();
 FILLCELL_X32 FILLER_155_97 ();
 FILLCELL_X32 FILLER_155_129 ();
 FILLCELL_X32 FILLER_155_161 ();
 FILLCELL_X16 FILLER_155_193 ();
 FILLCELL_X8 FILLER_155_209 ();
 FILLCELL_X2 FILLER_155_217 ();
 FILLCELL_X8 FILLER_155_271 ();
 FILLCELL_X2 FILLER_155_279 ();
 FILLCELL_X1 FILLER_155_281 ();
 FILLCELL_X8 FILLER_155_316 ();
 FILLCELL_X1 FILLER_155_324 ();
 FILLCELL_X2 FILLER_155_329 ();
 FILLCELL_X1 FILLER_155_379 ();
 FILLCELL_X32 FILLER_155_385 ();
 FILLCELL_X8 FILLER_155_417 ();
 FILLCELL_X4 FILLER_155_425 ();
 FILLCELL_X2 FILLER_155_429 ();
 FILLCELL_X4 FILLER_155_456 ();
 FILLCELL_X2 FILLER_155_476 ();
 FILLCELL_X1 FILLER_155_485 ();
 FILLCELL_X8 FILLER_155_489 ();
 FILLCELL_X1 FILLER_155_497 ();
 FILLCELL_X4 FILLER_155_502 ();
 FILLCELL_X8 FILLER_155_509 ();
 FILLCELL_X1 FILLER_155_517 ();
 FILLCELL_X1 FILLER_155_526 ();
 FILLCELL_X4 FILLER_155_536 ();
 FILLCELL_X2 FILLER_155_540 ();
 FILLCELL_X2 FILLER_155_570 ();
 FILLCELL_X1 FILLER_155_572 ();
 FILLCELL_X32 FILLER_155_612 ();
 FILLCELL_X32 FILLER_155_644 ();
 FILLCELL_X1 FILLER_155_676 ();
 FILLCELL_X1 FILLER_155_738 ();
 FILLCELL_X1 FILLER_155_764 ();
 FILLCELL_X1 FILLER_155_783 ();
 FILLCELL_X2 FILLER_155_788 ();
 FILLCELL_X1 FILLER_155_809 ();
 FILLCELL_X4 FILLER_155_817 ();
 FILLCELL_X2 FILLER_155_821 ();
 FILLCELL_X1 FILLER_155_823 ();
 FILLCELL_X1 FILLER_155_829 ();
 FILLCELL_X4 FILLER_155_864 ();
 FILLCELL_X1 FILLER_155_868 ();
 FILLCELL_X32 FILLER_155_876 ();
 FILLCELL_X32 FILLER_155_908 ();
 FILLCELL_X32 FILLER_155_940 ();
 FILLCELL_X32 FILLER_155_972 ();
 FILLCELL_X32 FILLER_155_1004 ();
 FILLCELL_X32 FILLER_155_1036 ();
 FILLCELL_X32 FILLER_155_1068 ();
 FILLCELL_X32 FILLER_155_1100 ();
 FILLCELL_X32 FILLER_155_1132 ();
 FILLCELL_X32 FILLER_155_1164 ();
 FILLCELL_X8 FILLER_155_1196 ();
 FILLCELL_X4 FILLER_155_1204 ();
 FILLCELL_X1 FILLER_155_1208 ();
 FILLCELL_X32 FILLER_156_1 ();
 FILLCELL_X32 FILLER_156_33 ();
 FILLCELL_X32 FILLER_156_65 ();
 FILLCELL_X32 FILLER_156_97 ();
 FILLCELL_X32 FILLER_156_129 ();
 FILLCELL_X32 FILLER_156_161 ();
 FILLCELL_X32 FILLER_156_193 ();
 FILLCELL_X8 FILLER_156_225 ();
 FILLCELL_X2 FILLER_156_233 ();
 FILLCELL_X1 FILLER_156_249 ();
 FILLCELL_X1 FILLER_156_275 ();
 FILLCELL_X4 FILLER_156_281 ();
 FILLCELL_X1 FILLER_156_285 ();
 FILLCELL_X4 FILLER_156_295 ();
 FILLCELL_X2 FILLER_156_299 ();
 FILLCELL_X1 FILLER_156_301 ();
 FILLCELL_X2 FILLER_156_307 ();
 FILLCELL_X4 FILLER_156_325 ();
 FILLCELL_X2 FILLER_156_329 ();
 FILLCELL_X1 FILLER_156_331 ();
 FILLCELL_X4 FILLER_156_334 ();
 FILLCELL_X2 FILLER_156_338 ();
 FILLCELL_X1 FILLER_156_340 ();
 FILLCELL_X32 FILLER_156_385 ();
 FILLCELL_X32 FILLER_156_417 ();
 FILLCELL_X4 FILLER_156_449 ();
 FILLCELL_X1 FILLER_156_482 ();
 FILLCELL_X4 FILLER_156_486 ();
 FILLCELL_X2 FILLER_156_490 ();
 FILLCELL_X1 FILLER_156_492 ();
 FILLCELL_X8 FILLER_156_496 ();
 FILLCELL_X2 FILLER_156_504 ();
 FILLCELL_X1 FILLER_156_510 ();
 FILLCELL_X8 FILLER_156_518 ();
 FILLCELL_X4 FILLER_156_537 ();
 FILLCELL_X2 FILLER_156_541 ();
 FILLCELL_X2 FILLER_156_550 ();
 FILLCELL_X2 FILLER_156_600 ();
 FILLCELL_X8 FILLER_156_616 ();
 FILLCELL_X4 FILLER_156_624 ();
 FILLCELL_X2 FILLER_156_628 ();
 FILLCELL_X1 FILLER_156_630 ();
 FILLCELL_X32 FILLER_156_632 ();
 FILLCELL_X16 FILLER_156_664 ();
 FILLCELL_X8 FILLER_156_680 ();
 FILLCELL_X2 FILLER_156_688 ();
 FILLCELL_X4 FILLER_156_694 ();
 FILLCELL_X2 FILLER_156_698 ();
 FILLCELL_X1 FILLER_156_700 ();
 FILLCELL_X1 FILLER_156_718 ();
 FILLCELL_X4 FILLER_156_768 ();
 FILLCELL_X2 FILLER_156_772 ();
 FILLCELL_X2 FILLER_156_788 ();
 FILLCELL_X1 FILLER_156_790 ();
 FILLCELL_X4 FILLER_156_813 ();
 FILLCELL_X4 FILLER_156_831 ();
 FILLCELL_X1 FILLER_156_835 ();
 FILLCELL_X1 FILLER_156_847 ();
 FILLCELL_X32 FILLER_156_855 ();
 FILLCELL_X32 FILLER_156_887 ();
 FILLCELL_X32 FILLER_156_919 ();
 FILLCELL_X32 FILLER_156_951 ();
 FILLCELL_X32 FILLER_156_983 ();
 FILLCELL_X32 FILLER_156_1015 ();
 FILLCELL_X32 FILLER_156_1047 ();
 FILLCELL_X32 FILLER_156_1079 ();
 FILLCELL_X32 FILLER_156_1111 ();
 FILLCELL_X32 FILLER_156_1143 ();
 FILLCELL_X32 FILLER_156_1175 ();
 FILLCELL_X2 FILLER_156_1207 ();
 FILLCELL_X32 FILLER_157_1 ();
 FILLCELL_X32 FILLER_157_33 ();
 FILLCELL_X32 FILLER_157_65 ();
 FILLCELL_X32 FILLER_157_97 ();
 FILLCELL_X32 FILLER_157_129 ();
 FILLCELL_X32 FILLER_157_161 ();
 FILLCELL_X32 FILLER_157_193 ();
 FILLCELL_X8 FILLER_157_225 ();
 FILLCELL_X4 FILLER_157_233 ();
 FILLCELL_X2 FILLER_157_247 ();
 FILLCELL_X2 FILLER_157_253 ();
 FILLCELL_X4 FILLER_157_272 ();
 FILLCELL_X2 FILLER_157_276 ();
 FILLCELL_X1 FILLER_157_296 ();
 FILLCELL_X4 FILLER_157_311 ();
 FILLCELL_X2 FILLER_157_315 ();
 FILLCELL_X1 FILLER_157_317 ();
 FILLCELL_X2 FILLER_157_327 ();
 FILLCELL_X1 FILLER_157_329 ();
 FILLCELL_X2 FILLER_157_334 ();
 FILLCELL_X1 FILLER_157_351 ();
 FILLCELL_X4 FILLER_157_367 ();
 FILLCELL_X2 FILLER_157_371 ();
 FILLCELL_X32 FILLER_157_380 ();
 FILLCELL_X32 FILLER_157_412 ();
 FILLCELL_X8 FILLER_157_444 ();
 FILLCELL_X2 FILLER_157_474 ();
 FILLCELL_X1 FILLER_157_485 ();
 FILLCELL_X1 FILLER_157_499 ();
 FILLCELL_X1 FILLER_157_504 ();
 FILLCELL_X1 FILLER_157_515 ();
 FILLCELL_X4 FILLER_157_531 ();
 FILLCELL_X2 FILLER_157_535 ();
 FILLCELL_X1 FILLER_157_544 ();
 FILLCELL_X1 FILLER_157_555 ();
 FILLCELL_X1 FILLER_157_560 ();
 FILLCELL_X4 FILLER_157_572 ();
 FILLCELL_X32 FILLER_157_611 ();
 FILLCELL_X32 FILLER_157_643 ();
 FILLCELL_X32 FILLER_157_675 ();
 FILLCELL_X2 FILLER_157_707 ();
 FILLCELL_X2 FILLER_157_738 ();
 FILLCELL_X8 FILLER_157_765 ();
 FILLCELL_X1 FILLER_157_773 ();
 FILLCELL_X2 FILLER_157_787 ();
 FILLCELL_X32 FILLER_157_799 ();
 FILLCELL_X32 FILLER_157_831 ();
 FILLCELL_X32 FILLER_157_863 ();
 FILLCELL_X32 FILLER_157_895 ();
 FILLCELL_X32 FILLER_157_927 ();
 FILLCELL_X32 FILLER_157_959 ();
 FILLCELL_X32 FILLER_157_991 ();
 FILLCELL_X32 FILLER_157_1023 ();
 FILLCELL_X32 FILLER_157_1055 ();
 FILLCELL_X32 FILLER_157_1087 ();
 FILLCELL_X32 FILLER_157_1119 ();
 FILLCELL_X32 FILLER_157_1151 ();
 FILLCELL_X16 FILLER_157_1183 ();
 FILLCELL_X8 FILLER_157_1199 ();
 FILLCELL_X2 FILLER_157_1207 ();
 FILLCELL_X32 FILLER_158_1 ();
 FILLCELL_X32 FILLER_158_33 ();
 FILLCELL_X32 FILLER_158_65 ();
 FILLCELL_X32 FILLER_158_97 ();
 FILLCELL_X32 FILLER_158_129 ();
 FILLCELL_X32 FILLER_158_161 ();
 FILLCELL_X32 FILLER_158_193 ();
 FILLCELL_X16 FILLER_158_225 ();
 FILLCELL_X4 FILLER_158_241 ();
 FILLCELL_X2 FILLER_158_262 ();
 FILLCELL_X1 FILLER_158_264 ();
 FILLCELL_X4 FILLER_158_273 ();
 FILLCELL_X1 FILLER_158_281 ();
 FILLCELL_X8 FILLER_158_291 ();
 FILLCELL_X1 FILLER_158_299 ();
 FILLCELL_X4 FILLER_158_304 ();
 FILLCELL_X1 FILLER_158_308 ();
 FILLCELL_X2 FILLER_158_317 ();
 FILLCELL_X1 FILLER_158_319 ();
 FILLCELL_X4 FILLER_158_324 ();
 FILLCELL_X1 FILLER_158_328 ();
 FILLCELL_X4 FILLER_158_333 ();
 FILLCELL_X32 FILLER_158_354 ();
 FILLCELL_X32 FILLER_158_386 ();
 FILLCELL_X32 FILLER_158_418 ();
 FILLCELL_X16 FILLER_158_450 ();
 FILLCELL_X4 FILLER_158_466 ();
 FILLCELL_X1 FILLER_158_470 ();
 FILLCELL_X1 FILLER_158_484 ();
 FILLCELL_X2 FILLER_158_540 ();
 FILLCELL_X2 FILLER_158_549 ();
 FILLCELL_X2 FILLER_158_561 ();
 FILLCELL_X1 FILLER_158_563 ();
 FILLCELL_X2 FILLER_158_571 ();
 FILLCELL_X1 FILLER_158_573 ();
 FILLCELL_X1 FILLER_158_584 ();
 FILLCELL_X1 FILLER_158_605 ();
 FILLCELL_X32 FILLER_158_632 ();
 FILLCELL_X32 FILLER_158_664 ();
 FILLCELL_X32 FILLER_158_696 ();
 FILLCELL_X32 FILLER_158_728 ();
 FILLCELL_X32 FILLER_158_760 ();
 FILLCELL_X32 FILLER_158_792 ();
 FILLCELL_X32 FILLER_158_824 ();
 FILLCELL_X32 FILLER_158_856 ();
 FILLCELL_X32 FILLER_158_888 ();
 FILLCELL_X32 FILLER_158_920 ();
 FILLCELL_X32 FILLER_158_952 ();
 FILLCELL_X32 FILLER_158_984 ();
 FILLCELL_X32 FILLER_158_1016 ();
 FILLCELL_X32 FILLER_158_1048 ();
 FILLCELL_X32 FILLER_158_1080 ();
 FILLCELL_X32 FILLER_158_1112 ();
 FILLCELL_X32 FILLER_158_1144 ();
 FILLCELL_X32 FILLER_158_1176 ();
 FILLCELL_X1 FILLER_158_1208 ();
 FILLCELL_X32 FILLER_159_1 ();
 FILLCELL_X32 FILLER_159_33 ();
 FILLCELL_X32 FILLER_159_65 ();
 FILLCELL_X32 FILLER_159_97 ();
 FILLCELL_X32 FILLER_159_129 ();
 FILLCELL_X32 FILLER_159_161 ();
 FILLCELL_X32 FILLER_159_193 ();
 FILLCELL_X32 FILLER_159_225 ();
 FILLCELL_X32 FILLER_159_257 ();
 FILLCELL_X32 FILLER_159_289 ();
 FILLCELL_X32 FILLER_159_321 ();
 FILLCELL_X32 FILLER_159_353 ();
 FILLCELL_X32 FILLER_159_385 ();
 FILLCELL_X32 FILLER_159_417 ();
 FILLCELL_X32 FILLER_159_449 ();
 FILLCELL_X2 FILLER_159_481 ();
 FILLCELL_X1 FILLER_159_483 ();
 FILLCELL_X2 FILLER_159_498 ();
 FILLCELL_X2 FILLER_159_510 ();
 FILLCELL_X16 FILLER_159_526 ();
 FILLCELL_X2 FILLER_159_542 ();
 FILLCELL_X1 FILLER_159_544 ();
 FILLCELL_X1 FILLER_159_555 ();
 FILLCELL_X2 FILLER_159_570 ();
 FILLCELL_X1 FILLER_159_599 ();
 FILLCELL_X32 FILLER_159_613 ();
 FILLCELL_X32 FILLER_159_645 ();
 FILLCELL_X32 FILLER_159_677 ();
 FILLCELL_X32 FILLER_159_709 ();
 FILLCELL_X32 FILLER_159_741 ();
 FILLCELL_X32 FILLER_159_773 ();
 FILLCELL_X32 FILLER_159_805 ();
 FILLCELL_X32 FILLER_159_837 ();
 FILLCELL_X32 FILLER_159_869 ();
 FILLCELL_X32 FILLER_159_901 ();
 FILLCELL_X32 FILLER_159_933 ();
 FILLCELL_X32 FILLER_159_965 ();
 FILLCELL_X32 FILLER_159_997 ();
 FILLCELL_X32 FILLER_159_1029 ();
 FILLCELL_X32 FILLER_159_1061 ();
 FILLCELL_X32 FILLER_159_1093 ();
 FILLCELL_X32 FILLER_159_1125 ();
 FILLCELL_X32 FILLER_159_1157 ();
 FILLCELL_X16 FILLER_159_1189 ();
 FILLCELL_X4 FILLER_159_1205 ();
 FILLCELL_X32 FILLER_160_1 ();
 FILLCELL_X32 FILLER_160_33 ();
 FILLCELL_X32 FILLER_160_65 ();
 FILLCELL_X32 FILLER_160_97 ();
 FILLCELL_X32 FILLER_160_129 ();
 FILLCELL_X32 FILLER_160_161 ();
 FILLCELL_X32 FILLER_160_193 ();
 FILLCELL_X32 FILLER_160_225 ();
 FILLCELL_X32 FILLER_160_257 ();
 FILLCELL_X32 FILLER_160_289 ();
 FILLCELL_X32 FILLER_160_321 ();
 FILLCELL_X32 FILLER_160_353 ();
 FILLCELL_X32 FILLER_160_385 ();
 FILLCELL_X32 FILLER_160_417 ();
 FILLCELL_X32 FILLER_160_449 ();
 FILLCELL_X16 FILLER_160_481 ();
 FILLCELL_X8 FILLER_160_497 ();
 FILLCELL_X4 FILLER_160_505 ();
 FILLCELL_X2 FILLER_160_509 ();
 FILLCELL_X1 FILLER_160_511 ();
 FILLCELL_X4 FILLER_160_547 ();
 FILLCELL_X1 FILLER_160_551 ();
 FILLCELL_X4 FILLER_160_561 ();
 FILLCELL_X1 FILLER_160_565 ();
 FILLCELL_X16 FILLER_160_602 ();
 FILLCELL_X8 FILLER_160_618 ();
 FILLCELL_X4 FILLER_160_626 ();
 FILLCELL_X1 FILLER_160_630 ();
 FILLCELL_X32 FILLER_160_632 ();
 FILLCELL_X32 FILLER_160_664 ();
 FILLCELL_X32 FILLER_160_696 ();
 FILLCELL_X32 FILLER_160_728 ();
 FILLCELL_X32 FILLER_160_760 ();
 FILLCELL_X32 FILLER_160_792 ();
 FILLCELL_X32 FILLER_160_824 ();
 FILLCELL_X32 FILLER_160_856 ();
 FILLCELL_X32 FILLER_160_888 ();
 FILLCELL_X32 FILLER_160_920 ();
 FILLCELL_X32 FILLER_160_952 ();
 FILLCELL_X32 FILLER_160_984 ();
 FILLCELL_X32 FILLER_160_1016 ();
 FILLCELL_X32 FILLER_160_1048 ();
 FILLCELL_X32 FILLER_160_1080 ();
 FILLCELL_X32 FILLER_160_1112 ();
 FILLCELL_X32 FILLER_160_1144 ();
 FILLCELL_X32 FILLER_160_1176 ();
 FILLCELL_X1 FILLER_160_1208 ();
 FILLCELL_X32 FILLER_161_1 ();
 FILLCELL_X32 FILLER_161_33 ();
 FILLCELL_X32 FILLER_161_65 ();
 FILLCELL_X32 FILLER_161_97 ();
 FILLCELL_X32 FILLER_161_129 ();
 FILLCELL_X32 FILLER_161_161 ();
 FILLCELL_X32 FILLER_161_193 ();
 FILLCELL_X32 FILLER_161_225 ();
 FILLCELL_X32 FILLER_161_257 ();
 FILLCELL_X32 FILLER_161_289 ();
 FILLCELL_X32 FILLER_161_321 ();
 FILLCELL_X32 FILLER_161_353 ();
 FILLCELL_X32 FILLER_161_385 ();
 FILLCELL_X32 FILLER_161_417 ();
 FILLCELL_X32 FILLER_161_449 ();
 FILLCELL_X8 FILLER_161_481 ();
 FILLCELL_X4 FILLER_161_489 ();
 FILLCELL_X1 FILLER_161_493 ();
 FILLCELL_X16 FILLER_161_511 ();
 FILLCELL_X2 FILLER_161_527 ();
 FILLCELL_X1 FILLER_161_529 ();
 FILLCELL_X4 FILLER_161_537 ();
 FILLCELL_X2 FILLER_161_541 ();
 FILLCELL_X4 FILLER_161_550 ();
 FILLCELL_X1 FILLER_161_554 ();
 FILLCELL_X8 FILLER_161_569 ();
 FILLCELL_X4 FILLER_161_577 ();
 FILLCELL_X2 FILLER_161_581 ();
 FILLCELL_X32 FILLER_161_600 ();
 FILLCELL_X32 FILLER_161_632 ();
 FILLCELL_X4 FILLER_161_664 ();
 FILLCELL_X4 FILLER_161_671 ();
 FILLCELL_X1 FILLER_161_675 ();
 FILLCELL_X2 FILLER_161_679 ();
 FILLCELL_X1 FILLER_161_681 ();
 FILLCELL_X32 FILLER_161_685 ();
 FILLCELL_X32 FILLER_161_717 ();
 FILLCELL_X32 FILLER_161_749 ();
 FILLCELL_X32 FILLER_161_781 ();
 FILLCELL_X32 FILLER_161_813 ();
 FILLCELL_X32 FILLER_161_845 ();
 FILLCELL_X32 FILLER_161_877 ();
 FILLCELL_X32 FILLER_161_909 ();
 FILLCELL_X32 FILLER_161_941 ();
 FILLCELL_X32 FILLER_161_973 ();
 FILLCELL_X32 FILLER_161_1005 ();
 FILLCELL_X32 FILLER_161_1037 ();
 FILLCELL_X32 FILLER_161_1069 ();
 FILLCELL_X32 FILLER_161_1101 ();
 FILLCELL_X32 FILLER_161_1133 ();
 FILLCELL_X32 FILLER_161_1165 ();
 FILLCELL_X8 FILLER_161_1197 ();
 FILLCELL_X4 FILLER_161_1205 ();
 FILLCELL_X32 FILLER_162_1 ();
 FILLCELL_X32 FILLER_162_33 ();
 FILLCELL_X32 FILLER_162_65 ();
 FILLCELL_X32 FILLER_162_97 ();
 FILLCELL_X32 FILLER_162_129 ();
 FILLCELL_X32 FILLER_162_161 ();
 FILLCELL_X32 FILLER_162_193 ();
 FILLCELL_X32 FILLER_162_225 ();
 FILLCELL_X32 FILLER_162_257 ();
 FILLCELL_X32 FILLER_162_289 ();
 FILLCELL_X32 FILLER_162_321 ();
 FILLCELL_X32 FILLER_162_353 ();
 FILLCELL_X32 FILLER_162_385 ();
 FILLCELL_X32 FILLER_162_417 ();
 FILLCELL_X32 FILLER_162_449 ();
 FILLCELL_X16 FILLER_162_481 ();
 FILLCELL_X8 FILLER_162_497 ();
 FILLCELL_X4 FILLER_162_505 ();
 FILLCELL_X1 FILLER_162_509 ();
 FILLCELL_X8 FILLER_162_513 ();
 FILLCELL_X2 FILLER_162_521 ();
 FILLCELL_X2 FILLER_162_540 ();
 FILLCELL_X1 FILLER_162_542 ();
 FILLCELL_X2 FILLER_162_556 ();
 FILLCELL_X1 FILLER_162_558 ();
 FILLCELL_X32 FILLER_162_566 ();
 FILLCELL_X32 FILLER_162_598 ();
 FILLCELL_X1 FILLER_162_630 ();
 FILLCELL_X2 FILLER_162_632 ();
 FILLCELL_X1 FILLER_162_634 ();
 FILLCELL_X8 FILLER_162_638 ();
 FILLCELL_X1 FILLER_162_646 ();
 FILLCELL_X2 FILLER_162_657 ();
 FILLCELL_X1 FILLER_162_659 ();
 FILLCELL_X8 FILLER_162_663 ();
 FILLCELL_X1 FILLER_162_675 ();
 FILLCELL_X4 FILLER_162_680 ();
 FILLCELL_X2 FILLER_162_687 ();
 FILLCELL_X4 FILLER_162_692 ();
 FILLCELL_X2 FILLER_162_696 ();
 FILLCELL_X4 FILLER_162_711 ();
 FILLCELL_X1 FILLER_162_715 ();
 FILLCELL_X32 FILLER_162_723 ();
 FILLCELL_X4 FILLER_162_755 ();
 FILLCELL_X2 FILLER_162_759 ();
 FILLCELL_X32 FILLER_162_764 ();
 FILLCELL_X32 FILLER_162_796 ();
 FILLCELL_X32 FILLER_162_828 ();
 FILLCELL_X32 FILLER_162_860 ();
 FILLCELL_X32 FILLER_162_892 ();
 FILLCELL_X32 FILLER_162_924 ();
 FILLCELL_X32 FILLER_162_956 ();
 FILLCELL_X32 FILLER_162_988 ();
 FILLCELL_X32 FILLER_162_1020 ();
 FILLCELL_X32 FILLER_162_1052 ();
 FILLCELL_X32 FILLER_162_1084 ();
 FILLCELL_X32 FILLER_162_1116 ();
 FILLCELL_X32 FILLER_162_1148 ();
 FILLCELL_X16 FILLER_162_1180 ();
 FILLCELL_X8 FILLER_162_1196 ();
 FILLCELL_X4 FILLER_162_1204 ();
 FILLCELL_X1 FILLER_162_1208 ();
 FILLCELL_X32 FILLER_163_1 ();
 FILLCELL_X32 FILLER_163_33 ();
 FILLCELL_X32 FILLER_163_65 ();
 FILLCELL_X32 FILLER_163_97 ();
 FILLCELL_X32 FILLER_163_129 ();
 FILLCELL_X32 FILLER_163_161 ();
 FILLCELL_X32 FILLER_163_193 ();
 FILLCELL_X32 FILLER_163_225 ();
 FILLCELL_X32 FILLER_163_257 ();
 FILLCELL_X32 FILLER_163_289 ();
 FILLCELL_X32 FILLER_163_321 ();
 FILLCELL_X32 FILLER_163_353 ();
 FILLCELL_X32 FILLER_163_385 ();
 FILLCELL_X32 FILLER_163_417 ();
 FILLCELL_X32 FILLER_163_449 ();
 FILLCELL_X16 FILLER_163_481 ();
 FILLCELL_X4 FILLER_163_497 ();
 FILLCELL_X1 FILLER_163_501 ();
 FILLCELL_X32 FILLER_163_505 ();
 FILLCELL_X8 FILLER_163_537 ();
 FILLCELL_X4 FILLER_163_545 ();
 FILLCELL_X4 FILLER_163_556 ();
 FILLCELL_X2 FILLER_163_560 ();
 FILLCELL_X1 FILLER_163_562 ();
 FILLCELL_X8 FILLER_163_566 ();
 FILLCELL_X2 FILLER_163_574 ();
 FILLCELL_X1 FILLER_163_580 ();
 FILLCELL_X4 FILLER_163_588 ();
 FILLCELL_X2 FILLER_163_592 ();
 FILLCELL_X1 FILLER_163_594 ();
 FILLCELL_X2 FILLER_163_607 ();
 FILLCELL_X1 FILLER_163_632 ();
 FILLCELL_X1 FILLER_163_654 ();
 FILLCELL_X4 FILLER_163_658 ();
 FILLCELL_X2 FILLER_163_662 ();
 FILLCELL_X1 FILLER_163_681 ();
 FILLCELL_X1 FILLER_163_702 ();
 FILLCELL_X2 FILLER_163_706 ();
 FILLCELL_X4 FILLER_163_720 ();
 FILLCELL_X8 FILLER_163_731 ();
 FILLCELL_X1 FILLER_163_739 ();
 FILLCELL_X4 FILLER_163_743 ();
 FILLCELL_X2 FILLER_163_747 ();
 FILLCELL_X1 FILLER_163_749 ();
 FILLCELL_X32 FILLER_163_756 ();
 FILLCELL_X2 FILLER_163_788 ();
 FILLCELL_X1 FILLER_163_790 ();
 FILLCELL_X4 FILLER_163_794 ();
 FILLCELL_X1 FILLER_163_798 ();
 FILLCELL_X8 FILLER_163_802 ();
 FILLCELL_X1 FILLER_163_810 ();
 FILLCELL_X32 FILLER_163_817 ();
 FILLCELL_X32 FILLER_163_849 ();
 FILLCELL_X32 FILLER_163_881 ();
 FILLCELL_X32 FILLER_163_913 ();
 FILLCELL_X32 FILLER_163_945 ();
 FILLCELL_X32 FILLER_163_977 ();
 FILLCELL_X32 FILLER_163_1009 ();
 FILLCELL_X32 FILLER_163_1041 ();
 FILLCELL_X32 FILLER_163_1073 ();
 FILLCELL_X32 FILLER_163_1105 ();
 FILLCELL_X32 FILLER_163_1137 ();
 FILLCELL_X32 FILLER_163_1169 ();
 FILLCELL_X8 FILLER_163_1201 ();
endmodule
